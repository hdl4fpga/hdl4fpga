library ieee;
use ieee.std_logic_1164.all;

package cgafonts4 is

	constant psf1cp850x8x16_80_to_FF : std_logic_vector(0 to 16*32*16-1) := (

		-- x"80" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"01100110" &
		B"11000010" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000010" &
		B"01100110" &
		B"00111100" &
		B"00011000" &
		B"01110000" &
		B"00000000" &
		B"00000000" &

		-- x"81" --
		B"00000000" &
		B"00000000" &
		B"11001100" &
		B"00000000" &
		B"00000000" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"82" --
		B"00000000" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"83" --
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"00000000" &
		B"01111000" &
		B"00001100" &
		B"01111100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"84" --
		B"00000000" &
		B"00000000" &
		B"11001100" &
		B"00000000" &
		B"00000000" &
		B"01111000" &
		B"00001100" &
		B"01111100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"85" --
		B"00000000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"01111000" &
		B"00001100" &
		B"01111100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"86" --
		B"00000000" &
		B"00111000" &
		B"01101100" &
		B"00111000" &
		B"00000000" &
		B"01111000" &
		B"00001100" &
		B"01111100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"87" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00011000" &
		B"01110000" &
		B"00000000" &
		B"00000000" &

		-- x"88" --
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"89" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"8a" --
		B"00000000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"8b" --
		B"00000000" &
		B"00000000" &
		B"01100110" &
		B"00000000" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"8c" --
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"01100110" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"8d" --
		B"00000000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"8e" --
		B"00000000" &
		B"11000110" &
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"8f" --
		B"00111000" &
		B"01101100" &
		B"00111000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"90" --
		B"00001100" &
		B"00011000" &
		B"00000000" &
		B"11111110" &
		B"01100110" &
		B"01100010" &
		B"01101000" &
		B"01111000" &
		B"01101000" &
		B"01100010" &
		B"01100110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"91" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11101100" &
		B"00110110" &
		B"00110110" &
		B"01111110" &
		B"11011000" &
		B"11011000" &
		B"01101110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"92" --
		B"00000000" &
		B"00000000" &
		B"00111110" &
		B"01101100" &
		B"11001100" &
		B"11001100" &
		B"11111110" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"93" --
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"94" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"95" --
		B"00000000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"96" --
		B"00000000" &
		B"00110000" &
		B"01111000" &
		B"11001100" &
		B"00000000" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"97" --
		B"00000000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"98" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"00001100" &
		B"01111000" &
		B"00000000" &

		-- x"99" --
		B"00000000" &
		B"11000110" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"9a" --
		B"00000000" &
		B"11000110" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"9b" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11001110" &
		B"11011110" &
		B"11110110" &
		B"11100110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"9c" --
		B"00000000" &
		B"00111000" &
		B"01101100" &
		B"01100100" &
		B"01100000" &
		B"11110000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"11100110" &
		B"11111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"9d" --
		B"00000000" &
		B"00000100" &
		B"01111100" &
		B"11001110" &
		B"11001110" &
		B"11010110" &
		B"11010110" &
		B"11010110" &
		B"11010110" &
		B"11100110" &
		B"11100110" &
		B"01111100" &
		B"01000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"9e" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"9f" --
		B"00000000" &
		B"00001110" &
		B"00011011" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11011000" &
		B"01110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a0" --
		B"00000000" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"00000000" &
		B"01111000" &
		B"00001100" &
		B"01111100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a1" --
		B"00000000" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a2" --
		B"00000000" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a3" --
		B"00000000" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"00000000" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a4" --
		B"00000000" &
		B"00000000" &
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"11011100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a5" --
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"11000110" &
		B"11100110" &
		B"11110110" &
		B"11111110" &
		B"11011110" &
		B"11001110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a6" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"01101100" &
		B"01101100" &
		B"00111110" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a7" --
		B"00000000" &
		B"00000000" &
		B"00111000" &
		B"01101100" &
		B"01101100" &
		B"00111000" &
		B"00000000" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a8" --
		B"00000000" &
		B"00000000" &
		B"00110000" &
		B"00110000" &
		B"00000000" &
		B"00110000" &
		B"00110000" &
		B"01100000" &
		B"11000000" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"a9" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"10000010" &
		B"10110010" &
		B"10101010" &
		B"10110010" &
		B"10101010" &
		B"10101010" &
		B"10000010" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"aa" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"ab" --
		B"00000000" &
		B"01100000" &
		B"11100000" &
		B"01100010" &
		B"01100110" &
		B"01101100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11011100" &
		B"10000110" &
		B"00001100" &
		B"00011000" &
		B"00111110" &
		B"00000000" &
		B"00000000" &

		-- x"ac" --
		B"00000000" &
		B"01100000" &
		B"11100000" &
		B"01100010" &
		B"01100110" &
		B"01101100" &
		B"00011000" &
		B"00110000" &
		B"01100110" &
		B"11001110" &
		B"10011010" &
		B"00111111" &
		B"00000110" &
		B"00000110" &
		B"00000000" &
		B"00000000" &

		-- x"ad" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00111100" &
		B"00111100" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"ae" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00110110" &
		B"01101100" &
		B"11011000" &
		B"01101100" &
		B"00110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"af" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11011000" &
		B"01101100" &
		B"00110110" &
		B"01101100" &
		B"11011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"b0" --
		B"00010001" &
		B"01000100" &
		B"00010001" &
		B"01000100" &
		B"00010001" &
		B"01000100" &
		B"00010001" &
		B"01000100" &
		B"00010001" &
		B"01000100" &
		B"00010001" &
		B"01000100" &
		B"00010001" &
		B"01000100" &
		B"00010001" &
		B"01000100" &

		-- x"b1" --
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &

		-- x"b2" --
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &

		-- x"b3" --
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		-- x"b4" --
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		-- x"b5" --
		B"01100000" &
		B"11000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"b6" --
		B"01111100" &
		B"11000110" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"b7" --
		B"00001100" &
		B"00000110" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"b8" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"10000010" &
		B"10011010" &
		B"10100010" &
		B"10100010" &
		B"10100010" &
		B"10011010" &
		B"10000010" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"b9" --
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"11110110" &
		B"00000110" &
		B"11110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		-- x"ba" --
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		-- x"bb" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"00000110" &
		B"11110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		-- x"bc" --
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"11110110" &
		B"00000110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"bd" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"be" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"bf" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		-- x"c0" --
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"c1" --
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"c2" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		-- x"c3" --
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		-- x"c4" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"c5" --
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11111111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		-- x"c6" --
		B"00000000" &
		B"00000000" &
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"01111000" &
		B"00001100" &
		B"01111100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"c7" --
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"c8" --
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110111" &
		B"00110000" &
		B"00111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"c9" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00111111" &
		B"00110000" &
		B"00110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		-- x"ca" --
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"11110111" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"cb" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"11110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		-- x"cc" --
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110111" &
		B"00110000" &
		B"00110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		-- x"cd" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"ce" --
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"11110111" &
		B"00000000" &
		B"11110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		-- x"cf" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d0" --
		B"00000000" &
		B"00000000" &
		B"00110100" &
		B"00011000" &
		B"00101100" &
		B"00000110" &
		B"00111110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d1" --
		B"00000000" &
		B"00000000" &
		B"11111000" &
		B"01101100" &
		B"01100110" &
		B"01100110" &
		B"11110110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01101100" &
		B"11111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d2" --
		B"00111000" &
		B"01101100" &
		B"00000000" &
		B"11111110" &
		B"01100110" &
		B"01100010" &
		B"01101000" &
		B"01111000" &
		B"01101000" &
		B"01100010" &
		B"01100110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d3" --
		B"00000000" &
		B"11000110" &
		B"00000000" &
		B"11111110" &
		B"01100110" &
		B"01100010" &
		B"01101000" &
		B"01111000" &
		B"01101000" &
		B"01100010" &
		B"01100110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d4" --
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"11111110" &
		B"01100110" &
		B"01100010" &
		B"01101000" &
		B"01111000" &
		B"01101000" &
		B"01100010" &
		B"01100110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d5" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d6" --
		B"00001100" &
		B"00011000" &
		B"00000000" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d7" --
		B"00111100" &
		B"01100110" &
		B"00000000" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d8" --
		B"00000000" &
		B"01100110" &
		B"00000000" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"d9" --
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"da" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		-- x"db" --
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &

		-- x"dc" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &

		-- x"dd" --
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"de" --
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"df" --
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"e0" --
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"e1" --
		B"00000000" &
		B"00000000" &
		B"01111000" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11011000" &
		B"11001100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11001100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"e2" --
		B"00111000" &
		B"01101100" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"e3" --
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"e4" --
		B"00000000" &
		B"00000000" &
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"e5" --
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"e6" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01100000" &
		B"01100000" &
		B"11000000" &
		B"00000000" &

		-- x"e7" --
		B"00000000" &
		B"00000000" &
		B"11100000" &
		B"01100000" &
		B"01100000" &
		B"01111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01100000" &
		B"01100000" &
		B"11110000" &
		B"00000000" &

		-- x"e8" --
		B"00000000" &
		B"00000000" &
		B"11110000" &
		B"01100000" &
		B"01111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01100000" &
		B"11110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"e9" --
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"ea" --
		B"00111000" &
		B"01101100" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"eb" --
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"ec" --
		B"00000000" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"00001100" &
		B"11111000" &
		B"00000000" &

		-- x"ed" --
		B"00001100" &
		B"00011000" &
		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"ee" --
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"ef" --
		B"00000000" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"f0" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"f1" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"f2" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"11111111" &
		B"00000000" &

		-- x"f3" --
		B"00000000" &
		B"11100000" &
		B"00110000" &
		B"01100010" &
		B"00110110" &
		B"11101100" &
		B"00011000" &
		B"00110000" &
		B"01100110" &
		B"11001110" &
		B"10011010" &
		B"00111111" &
		B"00000110" &
		B"00000110" &
		B"00000000" &
		B"00000000" &

		-- x"f4" --
		B"00000000" &
		B"00000000" &
		B"01111111" &
		B"11011011" &
		B"11011011" &
		B"11011011" &
		B"01111011" &
		B"00011011" &
		B"00011011" &
		B"00011011" &
		B"00011011" &
		B"00011011" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"f5" --
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"01100000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"00001100" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"f6" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"f7" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00001100" &
		B"01111000" &
		B"00000000" &
		B"00000000" &

		-- x"f8" --
		B"00000000" &
		B"00111000" &
		B"01101100" &
		B"01101100" &
		B"00111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"f9" --
		B"00000000" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"fa" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"fb" --
		B"00000000" &
		B"00011000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"fc" --
		B"00000000" &
		B"01111100" &
		B"00000110" &
		B"00111100" &
		B"00000110" &
		B"00000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"fd" --
		B"00000000" &
		B"00111100" &
		B"01100110" &
		B"00001100" &
		B"00011000" &
		B"00110010" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"fe" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"01111110" &
		B"01111110" &
		B"01111110" &
		B"01111110" &
		B"01111110" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"ff" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000"
		);

end;