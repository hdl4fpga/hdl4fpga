package test is
	constant std : natural := 0;
end;

