--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

library ieee;
use ieee.std_logic_1164.all;

package cgafonts is

--	constant psf1cp850x8x16 : std_logic_vector(0 to 256*8*16-1) := (
--		-- x"00" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"01" --
--		"00000000" &
--		"00000000" &
--		"01111110" &
--		"10000001" &
--		"10100101" &
--		"10000001" &
--		"10000001" &
--		"10111101" &
--		"10011001" &
--		"10000001" &
--		"10000001" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"02" --
--		"00000000" &
--		"00000000" &
--		"01111110" &
--		"11111111" &
--		"11011011" &
--		"11111111" &
--		"11111111" &
--		"11000011" &
--		"11100111" &
--		"11111111" &
--		"11111111" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"03" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01101100" &
--		"11111110" &
--		"11111110" &
--		"11111110" &
--		"11111110" &
--		"01111100" &
--		"00111000" &
--		"00010000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"04" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00010000" &
--		"00111000" &
--		"01111100" &
--		"11111110" &
--		"01111100" &
--		"00111000" &
--		"00010000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"05" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00111100" &
--		"00111100" &
--		"11100111" &
--		"11100111" &
--		"11100111" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"06" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00111100" &
--		"01111110" &
--		"11111111" &
--		"11111111" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"07" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00111100" &
--		"00111100" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"08" --
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11100111" &
--		"11000011" &
--		"11000011" &
--		"11100111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--
--		-- x"09" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"01100110" &
--		"01000010" &
--		"01000010" &
--		"01100110" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"0a" --
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11000011" &
--		"10011001" &
--		"10111101" &
--		"10111101" &
--		"10011001" &
--		"11000011" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--
--		-- x"0b" --
--		"00000000" &
--		"00000000" &
--		"00011110" &
--		"00001110" &
--		"00011010" &
--		"00110010" &
--		"01111000" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"0c" --
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"00111100" &
--		"00011000" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"0d" --
--		"00000000" &
--		"00000000" &
--		"00111111" &
--		"00110011" &
--		"00111111" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"01110000" &
--		"11110000" &
--		"11100000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"0e" --
--		"00000000" &
--		"00000000" &
--		"01111111" &
--		"01100011" &
--		"01111111" &
--		"01100011" &
--		"01100011" &
--		"01100011" &
--		"01100011" &
--		"01100111" &
--		"11100111" &
--		"11100110" &
--		"11000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"0f" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"11011011" &
--		"00111100" &
--		"11100111" &
--		"00111100" &
--		"11011011" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"10" --
--		"00000000" &
--		"10000000" &
--		"11000000" &
--		"11100000" &
--		"11110000" &
--		"11111000" &
--		"11111110" &
--		"11111000" &
--		"11110000" &
--		"11100000" &
--		"11000000" &
--		"10000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"11" --
--		"00000000" &
--		"00000010" &
--		"00000110" &
--		"00001110" &
--		"00011110" &
--		"00111110" &
--		"11111110" &
--		"00111110" &
--		"00011110" &
--		"00001110" &
--		"00000110" &
--		"00000010" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"12" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00111100" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"01111110" &
--		"00111100" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"13" --
--		"00000000" &
--		"00000000" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"00000000" &
--		"01100110" &
--		"01100110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"14" --
--		"00000000" &
--		"00000000" &
--		"01111111" &
--		"11011011" &
--		"11011011" &
--		"11011011" &
--		"01111011" &
--		"00011011" &
--		"00011011" &
--		"00011011" &
--		"00011011" &
--		"00011011" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"15" --
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"01100000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"01101100" &
--		"00111000" &
--		"00001100" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"16" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"11111110" &
--		"11111110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"17" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00111100" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"01111110" &
--		"00111100" &
--		"00011000" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"18" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00111100" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"19" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"01111110" &
--		"00111100" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"1a" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00001100" &
--		"11111110" &
--		"00001100" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"1b" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00110000" &
--		"01100000" &
--		"11111110" &
--		"01100000" &
--		"00110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"1c" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11000000" &
--		"11000000" &
--		"11000000" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"1d" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00101000" &
--		"01101100" &
--		"11111110" &
--		"01101100" &
--		"00101000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"1e" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00010000" &
--		"00111000" &
--		"00111000" &
--		"01111100" &
--		"01111100" &
--		"11111110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"1f" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"11111110" &
--		"01111100" &
--		"01111100" &
--		"00111000" &
--		"00111000" &
--		"00010000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"20" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"21" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00111100" &
--		"00111100" &
--		"00111100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"22" --
--		"00000000" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"00100100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"23" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01101100" &
--		"01101100" &
--		"11111110" &
--		"01101100" &
--		"01101100" &
--		"01101100" &
--		"11111110" &
--		"01101100" &
--		"01101100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"24" --
--		"00011000" &
--		"00011000" &
--		"01111100" &
--		"11000110" &
--		"11000010" &
--		"11000000" &
--		"01111100" &
--		"00000110" &
--		"00000110" &
--		"10000110" &
--		"11000110" &
--		"01111100" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"25" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11000010" &
--		"11000110" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"11000110" &
--		"10000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"26" --
--		"00000000" &
--		"00000000" &
--		"00111000" &
--		"01101100" &
--		"01101100" &
--		"00111000" &
--		"01110110" &
--		"11011100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"27" --
--		"00000000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"01100000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"28" --
--		"00000000" &
--		"00000000" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00011000" &
--		"00001100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"29" --
--		"00000000" &
--		"00000000" &
--		"00110000" &
--		"00011000" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"2a" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01100110" &
--		"00111100" &
--		"11111111" &
--		"00111100" &
--		"01100110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"2b" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"2c" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"2d" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"2e" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"2f" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000010" &
--		"00000110" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"11000000" &
--		"10000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"30" --
--		"00000000" &
--		"00000000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11010110" &
--		"11010110" &
--		"11000110" &
--		"11000110" &
--		"01101100" &
--		"00111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"31" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00111000" &
--		"01111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"32" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"00000110" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"11000000" &
--		"11000110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"33" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"00000110" &
--		"00000110" &
--		"00111100" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"34" --
--		"00000000" &
--		"00000000" &
--		"00001100" &
--		"00011100" &
--		"00111100" &
--		"01101100" &
--		"11001100" &
--		"11111110" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00011110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"35" --
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"11000000" &
--		"11000000" &
--		"11000000" &
--		"11111100" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"36" --
--		"00000000" &
--		"00000000" &
--		"00111000" &
--		"01100000" &
--		"11000000" &
--		"11000000" &
--		"11111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"37" --
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"11000110" &
--		"00000110" &
--		"00000110" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"38" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"39" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111110" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"00001100" &
--		"01111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"3a" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"3b" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"3c" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000110" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"00110000" &
--		"00011000" &
--		"00001100" &
--		"00000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"3d" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"3e" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01100000" &
--		"00110000" &
--		"00011000" &
--		"00001100" &
--		"00000110" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"3f" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"00001100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"40" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11011110" &
--		"11011110" &
--		"11011110" &
--		"11011100" &
--		"11000000" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"41" --
--		"00000000" &
--		"00000000" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"42" --
--		"00000000" &
--		"00000000" &
--		"11111100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01111100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"11111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"43" --
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"01100110" &
--		"11000010" &
--		"11000000" &
--		"11000000" &
--		"11000000" &
--		"11000000" &
--		"11000010" &
--		"01100110" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"44" --
--		"00000000" &
--		"00000000" &
--		"11111000" &
--		"01101100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01101100" &
--		"11111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"45" --
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"01100110" &
--		"01100010" &
--		"01101000" &
--		"01111000" &
--		"01101000" &
--		"01100000" &
--		"01100010" &
--		"01100110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"46" --
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"01100110" &
--		"01100010" &
--		"01101000" &
--		"01111000" &
--		"01101000" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"11110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"47" --
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"01100110" &
--		"11000010" &
--		"11000000" &
--		"11000000" &
--		"11011110" &
--		"11000110" &
--		"11000110" &
--		"01100110" &
--		"00111010" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"48" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"49" --
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"4a" --
--		"00000000" &
--		"00000000" &
--		"00011110" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"4b" --
--		"00000000" &
--		"00000000" &
--		"11100110" &
--		"01100110" &
--		"01100110" &
--		"01101100" &
--		"01111000" &
--		"01111000" &
--		"01101100" &
--		"01100110" &
--		"01100110" &
--		"11100110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"4c" --
--		"00000000" &
--		"00000000" &
--		"11110000" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"01100010" &
--		"01100110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"4d" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11101110" &
--		"11111110" &
--		"11111110" &
--		"11010110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"4e" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11100110" &
--		"11110110" &
--		"11111110" &
--		"11011110" &
--		"11001110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"4f" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"50" --
--		"00000000" &
--		"00000000" &
--		"11111100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01111100" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"11110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"51" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11010110" &
--		"11011110" &
--		"01111100" &
--		"00001100" &
--		"00001110" &
--		"00000000" &
--		"00000000" &
--
--		-- x"52" --
--		"00000000" &
--		"00000000" &
--		"11111100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01111100" &
--		"01101100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"11100110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"53" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"01100000" &
--		"00111000" &
--		"00001100" &
--		"00000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"54" --
--		"00000000" &
--		"00000000" &
--		"01111110" &
--		"01111110" &
--		"01011010" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"55" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"56" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01101100" &
--		"00111000" &
--		"00010000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"57" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11010110" &
--		"11010110" &
--		"11010110" &
--		"11111110" &
--		"11101110" &
--		"01101100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"58" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"01101100" &
--		"01111100" &
--		"00111000" &
--		"00111000" &
--		"01111100" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"59" --
--		"00000000" &
--		"00000000" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"00111100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"5a" --
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"11000110" &
--		"10000110" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"11000010" &
--		"11000110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"5b" --
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"5c" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"10000000" &
--		"11000000" &
--		"11100000" &
--		"01110000" &
--		"00111000" &
--		"00011100" &
--		"00001110" &
--		"00000110" &
--		"00000010" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"5d" --
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00001100" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"5e" --
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"5f" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111111" &
--		"00000000" &
--		"00000000" &
--
--		-- x"60" --
--		"00000000" &
--		"00110000" &
--		"00011000" &
--		"00001100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"61" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111000" &
--		"00001100" &
--		"01111100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"62" --
--		"00000000" &
--		"00000000" &
--		"11100000" &
--		"01100000" &
--		"01100000" &
--		"01111000" &
--		"01101100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"63" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000000" &
--		"11000000" &
--		"11000000" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"64" --
--		"00000000" &
--		"00000000" &
--		"00011100" &
--		"00001100" &
--		"00001100" &
--		"00111100" &
--		"01101100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"65" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11111110" &
--		"11000000" &
--		"11000000" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"66" --
--		"00000000" &
--		"00000000" &
--		"00011100" &
--		"00110110" &
--		"00110010" &
--		"00110000" &
--		"01111000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"01111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"67" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01110110" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01111100" &
--		"00001100" &
--		"11001100" &
--		"01111000" &
--		"00000000" &
--
--		-- x"68" --
--		"00000000" &
--		"00000000" &
--		"11100000" &
--		"01100000" &
--		"01100000" &
--		"01101100" &
--		"01110110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"11100110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"69" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"6a" --
--		"00000000" &
--		"00000000" &
--		"00000110" &
--		"00000110" &
--		"00000000" &
--		"00001110" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"01100110" &
--		"01100110" &
--		"00111100" &
--		"00000000" &
--
--		-- x"6b" --
--		"00000000" &
--		"00000000" &
--		"11100000" &
--		"01100000" &
--		"01100000" &
--		"01100110" &
--		"01101100" &
--		"01111000" &
--		"01111000" &
--		"01101100" &
--		"01100110" &
--		"11100110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"6c" --
--		"00000000" &
--		"00000000" &
--		"00111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"6d" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11101100" &
--		"11111110" &
--		"11010110" &
--		"11010110" &
--		"11010110" &
--		"11010110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"6e" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11011100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"6f" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"70" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11011100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01111100" &
--		"01100000" &
--		"01100000" &
--		"11110000" &
--		"00000000" &
--
--		-- x"71" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01110110" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01111100" &
--		"00001100" &
--		"00001100" &
--		"00011110" &
--		"00000000" &
--
--		-- x"72" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11011100" &
--		"01110110" &
--		"01100110" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"11110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"73" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"01100000" &
--		"00111000" &
--		"00001100" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"74" --
--		"00000000" &
--		"00000000" &
--		"00010000" &
--		"00110000" &
--		"00110000" &
--		"11111100" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110000" &
--		"00110110" &
--		"00011100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"75" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"76" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01101100" &
--		"00111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"77" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11010110" &
--		"11010110" &
--		"11010110" &
--		"11111110" &
--		"01101100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"78" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"01101100" &
--		"00111000" &
--		"00111000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"79" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111110" &
--		"00000110" &
--		"00001100" &
--		"11111000" &
--		"00000000" &
--
--		-- x"7a" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"11001100" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"11000110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"7b" --
--		"00000000" &
--		"00000000" &
--		"00001110" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"01110000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00001110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"7c" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"7d" --
--		"00000000" &
--		"00000000" &
--		"01110000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00001110" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"01110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"7e" --
--		"00000000" &
--		"01110110" &
--		"11011100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"7f" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"80" --
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"01100110" &
--		"11000010" &
--		"11000000" &
--		"11000000" &
--		"11000000" &
--		"11000000" &
--		"11000010" &
--		"01100110" &
--		"00111100" &
--		"00011000" &
--		"01110000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"81" --
--		"00000000" &
--		"00000000" &
--		"11001100" &
--		"00000000" &
--		"00000000" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"82" --
--		"00000000" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11111110" &
--		"11000000" &
--		"11000000" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"83" --
--		"00000000" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"00000000" &
--		"01111000" &
--		"00001100" &
--		"01111100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"84" --
--		"00000000" &
--		"00000000" &
--		"11001100" &
--		"00000000" &
--		"00000000" &
--		"01111000" &
--		"00001100" &
--		"01111100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"85" --
--		"00000000" &
--		"01100000" &
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"01111000" &
--		"00001100" &
--		"01111100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"86" --
--		"00000000" &
--		"00111000" &
--		"01101100" &
--		"00111000" &
--		"00000000" &
--		"01111000" &
--		"00001100" &
--		"01111100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"87" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000000" &
--		"11000000" &
--		"11000000" &
--		"11000110" &
--		"01111100" &
--		"00011000" &
--		"01110000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"88" --
--		"00000000" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11111110" &
--		"11000000" &
--		"11000000" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"89" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11111110" &
--		"11000000" &
--		"11000000" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"8a" --
--		"00000000" &
--		"01100000" &
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11111110" &
--		"11000000" &
--		"11000000" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"8b" --
--		"00000000" &
--		"00000000" &
--		"01100110" &
--		"00000000" &
--		"00000000" &
--		"00111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"8c" --
--		"00000000" &
--		"00011000" &
--		"00111100" &
--		"01100110" &
--		"00000000" &
--		"00111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"8d" --
--		"00000000" &
--		"01100000" &
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"00111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"8e" --
--		"00000000" &
--		"11000110" &
--		"00000000" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"8f" --
--		"00111000" &
--		"01101100" &
--		"00111000" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"90" --
--		"00001100" &
--		"00011000" &
--		"00000000" &
--		"11111110" &
--		"01100110" &
--		"01100010" &
--		"01101000" &
--		"01111000" &
--		"01101000" &
--		"01100010" &
--		"01100110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"91" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11101100" &
--		"00110110" &
--		"00110110" &
--		"01111110" &
--		"11011000" &
--		"11011000" &
--		"01101110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"92" --
--		"00000000" &
--		"00000000" &
--		"00111110" &
--		"01101100" &
--		"11001100" &
--		"11001100" &
--		"11111110" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"93" --
--		"00000000" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"94" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"95" --
--		"00000000" &
--		"01100000" &
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"96" --
--		"00000000" &
--		"00110000" &
--		"01111000" &
--		"11001100" &
--		"00000000" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"97" --
--		"00000000" &
--		"01100000" &
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"98" --
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111110" &
--		"00000110" &
--		"00001100" &
--		"01111000" &
--		"00000000" &
--
--		-- x"99" --
--		"00000000" &
--		"11000110" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"9a" --
--		"00000000" &
--		"11000110" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"9b" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"11001110" &
--		"11011110" &
--		"11110110" &
--		"11100110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"9c" --
--		"00000000" &
--		"00111000" &
--		"01101100" &
--		"01100100" &
--		"01100000" &
--		"11110000" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"01100000" &
--		"11100110" &
--		"11111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"9d" --
--		"00000000" &
--		"00000100" &
--		"01111100" &
--		"11001110" &
--		"11001110" &
--		"11010110" &
--		"11010110" &
--		"11010110" &
--		"11010110" &
--		"11100110" &
--		"11100110" &
--		"01111100" &
--		"01000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"9e" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"01101100" &
--		"00111000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"9f" --
--		"00000000" &
--		"00001110" &
--		"00011011" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"11011000" &
--		"01110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a0" --
--		"00000000" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"00000000" &
--		"01111000" &
--		"00001100" &
--		"01111100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a1" --
--		"00000000" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"00111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a2" --
--		"00000000" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a3" --
--		"00000000" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"00000000" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a4" --
--		"00000000" &
--		"00000000" &
--		"01110110" &
--		"11011100" &
--		"00000000" &
--		"11011100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a5" --
--		"01110110" &
--		"11011100" &
--		"00000000" &
--		"11000110" &
--		"11100110" &
--		"11110110" &
--		"11111110" &
--		"11011110" &
--		"11001110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a6" --
--		"00000000" &
--		"00000000" &
--		"00111100" &
--		"01101100" &
--		"01101100" &
--		"00111110" &
--		"00000000" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a7" --
--		"00000000" &
--		"00000000" &
--		"00111000" &
--		"01101100" &
--		"01101100" &
--		"00111000" &
--		"00000000" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a8" --
--		"00000000" &
--		"00000000" &
--		"00110000" &
--		"00110000" &
--		"00000000" &
--		"00110000" &
--		"00110000" &
--		"01100000" &
--		"11000000" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"a9" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"10000010" &
--		"10110010" &
--		"10101010" &
--		"10110010" &
--		"10101010" &
--		"10101010" &
--		"10000010" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"aa" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"00000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ab" --
--		"00000000" &
--		"01100000" &
--		"11100000" &
--		"01100010" &
--		"01100110" &
--		"01101100" &
--		"00011000" &
--		"00110000" &
--		"01100000" &
--		"11011100" &
--		"10000110" &
--		"00001100" &
--		"00011000" &
--		"00111110" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ac" --
--		"00000000" &
--		"01100000" &
--		"11100000" &
--		"01100010" &
--		"01100110" &
--		"01101100" &
--		"00011000" &
--		"00110000" &
--		"01100110" &
--		"11001110" &
--		"10011010" &
--		"00111111" &
--		"00000110" &
--		"00000110" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ad" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00111100" &
--		"00111100" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ae" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00110110" &
--		"01101100" &
--		"11011000" &
--		"01101100" &
--		"00110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"af" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11011000" &
--		"01101100" &
--		"00110110" &
--		"01101100" &
--		"11011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"b0" --
--		"00010001" &
--		"01000100" &
--		"00010001" &
--		"01000100" &
--		"00010001" &
--		"01000100" &
--		"00010001" &
--		"01000100" &
--		"00010001" &
--		"01000100" &
--		"00010001" &
--		"01000100" &
--		"00010001" &
--		"01000100" &
--		"00010001" &
--		"01000100" &
--
--		-- x"b1" --
--		"01010101" &
--		"10101010" &
--		"01010101" &
--		"10101010" &
--		"01010101" &
--		"10101010" &
--		"01010101" &
--		"10101010" &
--		"01010101" &
--		"10101010" &
--		"01010101" &
--		"10101010" &
--		"01010101" &
--		"10101010" &
--		"01010101" &
--		"10101010" &
--
--		-- x"b2" --
--		"11011101" &
--		"01110111" &
--		"11011101" &
--		"01110111" &
--		"11011101" &
--		"01110111" &
--		"11011101" &
--		"01110111" &
--		"11011101" &
--		"01110111" &
--		"11011101" &
--		"01110111" &
--		"11011101" &
--		"01110111" &
--		"11011101" &
--		"01110111" &
--
--		-- x"b3" --
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--
--		-- x"b4" --
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"11111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--
--		-- x"b5" --
--		"01100000" &
--		"11000000" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"b6" --
--		"01111100" &
--		"11000110" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"b7" --
--		"00001100" &
--		"00000110" &
--		"00010000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"b8" --
--		"00000000" &
--		"00000000" &
--		"01111100" &
--		"10000010" &
--		"10011010" &
--		"10100010" &
--		"10100010" &
--		"10100010" &
--		"10011010" &
--		"10000010" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"b9" --
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"11110110" &
--		"00000110" &
--		"11110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--
--		-- x"ba" --
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--
--		-- x"bb" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"00000110" &
--		"11110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--
--		-- x"bc" --
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"11110110" &
--		"00000110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"bd" --
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"01111100" &
--		"11000110" &
--		"11000000" &
--		"11000000" &
--		"11000110" &
--		"01111100" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"be" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01100110" &
--		"01100110" &
--		"00111100" &
--		"00011000" &
--		"01111110" &
--		"00011000" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"bf" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--
--		-- x"c0" --
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011111" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"c1" --
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"11111111" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"c2" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111111" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--
--		-- x"c3" --
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011111" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--
--		-- x"c4" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111111" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"c5" --
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"11111111" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--
--		-- x"c6" --
--		"00000000" &
--		"00000000" &
--		"01110110" &
--		"11011100" &
--		"00000000" &
--		"01111000" &
--		"00001100" &
--		"01111100" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"01110110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"c7" --
--		"01110110" &
--		"11011100" &
--		"00000000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"11111110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"c8" --
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110111" &
--		"00110000" &
--		"00111111" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"c9" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00111111" &
--		"00110000" &
--		"00110111" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--
--		-- x"ca" --
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"11110111" &
--		"00000000" &
--		"11111111" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"cb" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111111" &
--		"00000000" &
--		"11110111" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--
--		-- x"cc" --
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110111" &
--		"00110000" &
--		"00110111" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--
--		-- x"cd" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111111" &
--		"00000000" &
--		"11111111" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ce" --
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"11110111" &
--		"00000000" &
--		"11110111" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--		"00110110" &
--
--		-- x"cf" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11000110" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d0" --
--		"00000000" &
--		"00000000" &
--		"00110100" &
--		"00011000" &
--		"00101100" &
--		"00000110" &
--		"00111110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d1" --
--		"00000000" &
--		"00000000" &
--		"11111000" &
--		"01101100" &
--		"01100110" &
--		"01100110" &
--		"11110110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01101100" &
--		"11111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d2" --
--		"00111000" &
--		"01101100" &
--		"00000000" &
--		"11111110" &
--		"01100110" &
--		"01100010" &
--		"01101000" &
--		"01111000" &
--		"01101000" &
--		"01100010" &
--		"01100110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d3" --
--		"00000000" &
--		"11000110" &
--		"00000000" &
--		"11111110" &
--		"01100110" &
--		"01100010" &
--		"01101000" &
--		"01111000" &
--		"01101000" &
--		"01100010" &
--		"01100110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d4" --
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"11111110" &
--		"01100110" &
--		"01100010" &
--		"01101000" &
--		"01111000" &
--		"01101000" &
--		"01100010" &
--		"01100110" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d5" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d6" --
--		"00001100" &
--		"00011000" &
--		"00000000" &
--		"00111100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d7" --
--		"00111100" &
--		"01100110" &
--		"00000000" &
--		"00111100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d8" --
--		"00000000" &
--		"01100110" &
--		"00000000" &
--		"00111100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"d9" --
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"11111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"da" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011111" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--
--		-- x"db" --
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--
--		-- x"dc" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--
--		-- x"dd" --
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"de" --
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"00111100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"df" --
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"11111111" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"e0" --
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"e1" --
--		"00000000" &
--		"00000000" &
--		"01111000" &
--		"11001100" &
--		"11001100" &
--		"11001100" &
--		"11011000" &
--		"11001100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11001100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"e2" --
--		"00111000" &
--		"01101100" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"e3" --
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"e4" --
--		"00000000" &
--		"00000000" &
--		"01110110" &
--		"11011100" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"e5" --
--		"01110110" &
--		"11011100" &
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"e6" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01111100" &
--		"01100000" &
--		"01100000" &
--		"11000000" &
--		"00000000" &
--
--		-- x"e7" --
--		"00000000" &
--		"00000000" &
--		"11100000" &
--		"01100000" &
--		"01100000" &
--		"01111100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01111100" &
--		"01100000" &
--		"01100000" &
--		"11110000" &
--		"00000000" &
--
--		-- x"e8" --
--		"00000000" &
--		"00000000" &
--		"11110000" &
--		"01100000" &
--		"01111100" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01111100" &
--		"01100000" &
--		"11110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"e9" --
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ea" --
--		"00111000" &
--		"01101100" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"eb" --
--		"00110000" &
--		"00011000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ec" --
--		"00000000" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"11000110" &
--		"01111110" &
--		"00000110" &
--		"00001100" &
--		"11111000" &
--		"00000000" &
--
--		-- x"ed" --
--		"00001100" &
--		"00011000" &
--		"00000000" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"01100110" &
--		"00111100" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ee" --
--		"00000000" &
--		"11111111" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ef" --
--		"00000000" &
--		"00001100" &
--		"00011000" &
--		"00110000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f0" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f1" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00011000" &
--		"01111110" &
--		"00011000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f2" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"11111111" &
--		"00000000" &
--		"11111111" &
--		"00000000" &
--
--		-- x"f3" --
--		"00000000" &
--		"11100000" &
--		"00110000" &
--		"01100010" &
--		"00110110" &
--		"11101100" &
--		"00011000" &
--		"00110000" &
--		"01100110" &
--		"11001110" &
--		"10011010" &
--		"00111111" &
--		"00000110" &
--		"00000110" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f4" --
--		"00000000" &
--		"00000000" &
--		"01111111" &
--		"11011011" &
--		"11011011" &
--		"11011011" &
--		"01111011" &
--		"00011011" &
--		"00011011" &
--		"00011011" &
--		"00011011" &
--		"00011011" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f5" --
--		"00000000" &
--		"01111100" &
--		"11000110" &
--		"01100000" &
--		"00111000" &
--		"01101100" &
--		"11000110" &
--		"11000110" &
--		"01101100" &
--		"00111000" &
--		"00001100" &
--		"11000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f6" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00000000" &
--		"01111110" &
--		"00000000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f7" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00001100" &
--		"01111000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f8" --
--		"00000000" &
--		"00111000" &
--		"01101100" &
--		"01101100" &
--		"00111000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"f9" --
--		"00000000" &
--		"11000110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"fa" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00011000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"fb" --
--		"00000000" &
--		"00011000" &
--		"00111000" &
--		"00011000" &
--		"00011000" &
--		"00011000" &
--		"00111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"fc" --
--		"00000000" &
--		"01111100" &
--		"00000110" &
--		"00111100" &
--		"00000110" &
--		"00000110" &
--		"01111100" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"fd" --
--		"00000000" &
--		"00111100" &
--		"01100110" &
--		"00001100" &
--		"00011000" &
--		"00110010" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"fe" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"01111110" &
--		"01111110" &
--		"01111110" &
--		"01111110" &
--		"01111110" &
--		"01111110" &
--		"01111110" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--
--		-- x"ff" --
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000" &
--		"00000000");

	constant psf1digit8x8 : std_logic_vector(0 to 16*8*8-1) := (
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00011000" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00000000" &

		"01111100" &
		"11000110" &
		"00000110" &
		"01111100" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &

		"11111100" &
		"00000110" &
		"00000110" &
		"00111100" &
		"00000110" &
		"00000110" &
		"11111100" &
		"00000000" &

		"00001100" &
		"11001100" &
		"11001100" &
		"11001100" &
		"11111110" &
		"00001100" &
		"00001100" &
		"00000000" &

		"11111110" &
		"11000000" &
		"11111100" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"01111100" &
		"11000000" &
		"11000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111110" &
		"00000110" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"00110000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"00000110" &
		"01111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00111110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111111" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000");


	constant psf1cp850x8x8 : std_logic_vector(0 to 256*8*8-1) := (

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"01111110" &
		"10000001" &
		"10100101" &
		"10000001" &
		"10011101" &
		"10111001" &
		"10000001" &
		"01111110" &

		"01111110" &
		"11111111" &
		"11011011" &
		"11111111" &
		"11100011" &
		"11000111" &
		"11111111" &
		"01111110" &

		"01101100" &
		"11111110" &
		"11111110" &
		"11111110" &
		"01111100" &
		"00111000" &
		"00010000" &
		"00000000" &

		"00010000" &
		"00111000" &
		"01111100" &
		"11111110" &
		"01111100" &
		"00111000" &
		"00010000" &
		"00000000" &

		"00111000" &
		"01111100" &
		"00111000" &
		"11111110" &
		"11111110" &
		"00010000" &
		"00010000" &
		"01111100" &

		"00000000" &
		"00011000" &
		"00111100" &
		"01111110" &
		"11111111" &
		"01111110" &
		"00011000" &
		"01111110" &

		"00000000" &
		"00000000" &
		"00011000" &
		"00111100" &
		"00111100" &
		"00011000" &
		"00000000" &
		"00000000" &

		"11111111" &
		"11111111" &
		"11100111" &
		"11000011" &
		"11000011" &
		"11100111" &
		"11111111" &
		"11111111" &

		"00000000" &
		"00111100" &
		"01100110" &
		"01000010" &
		"01000010" &
		"01100110" &
		"00111100" &
		"00000000" &

		"11111111" &
		"11000011" &
		"10011001" &
		"10111101" &
		"10111101" &
		"10011001" &
		"11000011" &
		"11111111" &

		"00001111" &
		"00000111" &
		"00001111" &
		"01111101" &
		"11001100" &
		"11001100" &
		"11001100" &
		"01111000" &

		"00111100" &
		"01100110" &
		"01100110" &
		"01100110" &
		"00111100" &
		"00011000" &
		"01111110" &
		"00011000" &

		"00111111" &
		"00110011" &
		"00111111" &
		"00110000" &
		"00110000" &
		"01110000" &
		"11110000" &
		"11100000" &

		"01111111" &
		"01100011" &
		"01111111" &
		"01100011" &
		"01100011" &
		"01100111" &
		"11100110" &
		"11000000" &

		"10011001" &
		"01011010" &
		"00111100" &
		"11100111" &
		"11100111" &
		"00111100" &
		"01011010" &
		"10011001" &

		"10000000" &
		"11100000" &
		"11111000" &
		"11111110" &
		"11111000" &
		"11100000" &
		"10000000" &
		"00000000" &

		"00000010" &
		"00001110" &
		"00111110" &
		"11111110" &
		"00111110" &
		"00001110" &
		"00000010" &
		"00000000" &

		"00011000" &
		"00111100" &
		"01111110" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00111100" &
		"00011000" &

		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"00000000" &
		"01100110" &
		"00000000" &

		"01111111" &
		"11011011" &
		"11011011" &
		"01111011" &
		"00011011" &
		"00011011" &
		"00011011" &
		"00000000" &

		"00111111" &
		"01100000" &
		"01111100" &
		"01100110" &
		"01100110" &
		"00111110" &
		"00000110" &
		"11111100" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"01111110" &
		"01111110" &
		"01111110" &
		"00000000" &

		"00011000" &
		"00111100" &
		"01111110" &
		"00011000" &
		"01111110" &
		"00111100" &
		"00011000" &
		"11111111" &

		"00011000" &
		"00111100" &
		"01111110" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00111100" &
		"00011000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00001100" &
		"11111110" &
		"00001100" &
		"00011000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00110000" &
		"01100000" &
		"11111110" &
		"01100000" &
		"00110000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00100100" &
		"01100110" &
		"11111111" &
		"01100110" &
		"00100100" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00111100" &
		"01111110" &
		"11111111" &
		"11111111" &
		"00000000" &
		"00000000" &

		"00000000" &
		"11111111" &
		"11111111" &
		"01111110" &
		"00111100" &
		"00011000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00011000" &
		"00000000" &

		"01101100" &
		"01101100" &
		"01101100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"01101100" &
		"01101100" &
		"11111110" &
		"01101100" &
		"11111110" &
		"01101100" &
		"01101100" &
		"00000000" &

		"00011000" &
		"01111110" &
		"11000000" &
		"01111100" &
		"00000110" &
		"11111100" &
		"00011000" &
		"00000000" &

		"00000000" &
		"11000110" &
		"11001100" &
		"00011000" &
		"00110000" &
		"01100110" &
		"11000110" &
		"00000000" &

		"00111000" &
		"01101100" &
		"00111000" &
		"01110110" &
		"11011100" &
		"11001100" &
		"01110110" &
		"00000000" &

		"00110000" &
		"00110000" &
		"01100000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00001100" &
		"00011000" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00011000" &
		"00001100" &
		"00000000" &

		"00110000" &
		"00011000" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00011000" &
		"00110000" &
		"00000000" &

		"00000000" &
		"01100110" &
		"00111100" &
		"11111111" &
		"00111100" &
		"01100110" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00110000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"01111110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"01100000" &
		"11000000" &
		"10000000" &
		"00000000" &

		"01111100" &
		"11001110" &
		"11011110" &
		"11110110" &
		"11100110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00011000" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00000000" &

		"01111100" &
		"11000110" &
		"00000110" &
		"01111100" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &

		"11111100" &
		"00000110" &
		"00000110" &
		"00111100" &
		"00000110" &
		"00000110" &
		"11111100" &
		"00000000" &

		"00001100" &
		"11001100" &
		"11001100" &
		"11001100" &
		"11111110" &
		"00001100" &
		"00001100" &
		"00000000" &

		"11111110" &
		"11000000" &
		"11111100" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"01111100" &
		"11000000" &
		"11000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111110" &
		"00000110" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"00110000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"00000110" &
		"01111100" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00110000" &

		"00001100" &
		"00011000" &
		"00110000" &
		"01100000" &
		"00110000" &
		"00011000" &
		"00001100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"00000000" &
		"01111110" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00110000" &
		"00011000" &
		"00001100" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"00000000" &

		"00111100" &
		"01100110" &
		"00001100" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00011000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11011110" &
		"11011110" &
		"11011110" &
		"11000000" &
		"01111110" &
		"00000000" &

		"00111000" &
		"01101100" &
		"11000110" &
		"11000110" &
		"11111110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111000" &
		"11001100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11001100" &
		"11111000" &
		"00000000" &

		"11111110" &
		"11000000" &
		"11000000" &
		"11111000" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &

		"11111110" &
		"11000000" &
		"11000000" &
		"11111000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000000" &
		"11000000" &
		"11001110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"11111110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"01111110" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00000000" &

		"00000110" &
		"00000110" &
		"00000110" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11000110" &
		"11001100" &
		"11011000" &
		"11110000" &
		"11011000" &
		"11001100" &
		"11000110" &
		"00000000" &

		"11000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &

		"11000110" &
		"11101110" &
		"11111110" &
		"11111110" &
		"11010110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"11000110" &
		"11100110" &
		"11110110" &
		"11011110" &
		"11001110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"11000000" &
		"11000000" &
		"11000000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11010110" &
		"11011110" &
		"01111100" &
		"00000110" &

		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"11011000" &
		"11001100" &
		"11000110" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000000" &
		"01111100" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111111" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11111110" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00111000" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11010110" &
		"11111110" &
		"01101100" &
		"00000000" &

		"11000110" &
		"11000110" &
		"01101100" &
		"00111000" &
		"01101100" &
		"11000110" &
		"11000110" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00011000" &
		"00110000" &
		"11100000" &
		"00000000" &

		"11111110" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"01100000" &
		"11111110" &
		"00000000" &

		"00111100" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00111100" &
		"00000000" &

		"11000000" &
		"01100000" &
		"00110000" &
		"00011000" &
		"00001100" &
		"00000110" &
		"00000010" &
		"00000000" &

		"00111100" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00111100" &
		"00000000" &

		"00010000" &
		"00111000" &
		"01101100" &
		"11000110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111111" &

		"00011000" &
		"00011000" &
		"00001100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"00000110" &
		"01111110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"11000000" &
		"11000000" &
		"11000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000000" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00000110" &
		"00000110" &
		"00000110" &
		"01111110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11111110" &
		"11000000" &
		"01111100" &
		"00000000" &

		"00011100" &
		"00110110" &
		"00110000" &
		"01111000" &
		"00110000" &
		"00110000" &
		"01111000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"11111100" &

		"11000000" &
		"11000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"00011000" &
		"00000000" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00111100" &
		"00000000" &

		"00000110" &
		"00000000" &
		"00000110" &
		"00000110" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &

		"11000000" &
		"11000000" &
		"11001100" &
		"11011000" &
		"11111000" &
		"11001100" &
		"11000110" &
		"00000000" &

		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11001100" &
		"11111110" &
		"11111110" &
		"11010110" &
		"11010110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"11000000" &
		"11000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"00000110" &

		"00000000" &
		"00000000" &
		"11111100" &
		"11000110" &
		"11000000" &
		"11000000" &
		"11000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"11000000" &
		"01111100" &
		"00000110" &
		"11111100" &
		"00000000" &

		"00011000" &
		"00011000" &
		"01111110" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00001110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00111000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11010110" &
		"11111110" &
		"01101100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"01101100" &
		"00111000" &
		"01101100" &
		"11000110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"11111100" &

		"00000000" &
		"00000000" &
		"11111110" &
		"00001100" &
		"00111000" &
		"01100000" &
		"11111110" &
		"00000000" &

		"00001110" &
		"00011000" &
		"00011000" &
		"01110000" &
		"00011000" &
		"00011000" &
		"00001110" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"01110000" &
		"00011000" &
		"00011000" &
		"00001110" &
		"00011000" &
		"00011000" &
		"01110000" &
		"00000000" &

		"01110110" &
		"11011100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00010000" &
		"00111000" &
		"01101100" &
		"11000110" &
		"11000110" &
		"11111110" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11010110" &
		"01111100" &
		"00110000" &

		"11000110" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00001110" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11111110" &
		"11000000" &
		"01111100" &
		"00000000" &

		"01111110" &
		"10000001" &
		"00111100" &
		"00000110" &
		"01111110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"01100110" &
		"00000000" &
		"01111100" &
		"00000110" &
		"01111110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"11100000" &
		"00000000" &
		"01111100" &
		"00000110" &
		"01111110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00011000" &
		"00011000" &
		"01111100" &
		"00000110" &
		"01111110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000000" &
		"11010110" &
		"01111100" &
		"00110000" &

		"01111110" &
		"10000001" &
		"01111100" &
		"11000110" &
		"11111110" &
		"11000000" &
		"01111100" &
		"00000000" &

		"01100110" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11111110" &
		"11000000" &
		"01111100" &
		"00000000" &

		"11100000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11111110" &
		"11000000" &
		"01111100" &
		"00000000" &

		"01100110" &
		"00000000" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00111100" &
		"00000000" &

		"01111100" &
		"10000010" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00111100" &
		"00000000" &

		"01110000" &
		"00000000" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00111100" &
		"00000000" &

		"11000110" &
		"00010000" &
		"01111100" &
		"11000110" &
		"11111110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"00111000" &
		"00111000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11111110" &
		"11000110" &
		"00000000" &

		"00001110" &
		"00000000" &
		"11111110" &
		"11000000" &
		"11111000" &
		"11000000" &
		"11111110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111111" &
		"00001100" &
		"01111111" &
		"11001100" &
		"01111111" &
		"00000000" &

		"00111111" &
		"01101100" &
		"11001100" &
		"11111111" &
		"11001100" &
		"11001100" &
		"11001111" &
		"00000000" &

		"01111100" &
		"10000010" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"01100110" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11100000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"01111100" &
		"10000010" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"11100000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"01100110" &
		"00000000" &
		"01100110" &
		"01100110" &
		"01100110" &
		"00111110" &
		"00000110" &
		"01111100" &

		"11000110" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11000110" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11111110" &
		"00000000" &

		"00011000" &
		"00011000" &
		"01111110" &
		"11011000" &
		"11011000" &
		"11011000" &
		"01111110" &
		"00011000" &

		"00111000" &
		"01101100" &
		"01100000" &
		"11110000" &
		"01100000" &
		"01100110" &
		"11111100" &
		"00000000" &

		"01100110" &
		"01100110" &
		"00111100" &
		"00011000" &
		"01111110" &
		"00011000" &
		"01111110" &
		"00011000" &

		"11111000" &
		"11001100" &
		"11001100" &
		"11111010" &
		"11000110" &
		"11001111" &
		"11000110" &
		"11000011" &

		"00001110" &
		"00011011" &
		"00011000" &
		"00111100" &
		"00011000" &
		"00011000" &
		"11011000" &
		"01110000" &

		"00001110" &
		"00000000" &
		"01111100" &
		"00000110" &
		"01111110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00011100" &
		"00000000" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00111100" &
		"00000000" &

		"00001110" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00001110" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00000000" &
		"11111110" &
		"00000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"11111110" &
		"00000000" &
		"11000110" &
		"11100110" &
		"11110110" &
		"11011110" &
		"11001110" &
		"00000000" &

		"00111100" &
		"01101100" &
		"01101100" &
		"00111110" &
		"00000000" &
		"01111110" &
		"00000000" &
		"00000000" &

		"00111100" &
		"01100110" &
		"01100110" &
		"00111100" &
		"00000000" &
		"01111110" &
		"00000000" &
		"00000000" &

		"00011000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00110000" &
		"01100110" &
		"00111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"11111100" &
		"11000000" &
		"11000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"11111100" &
		"00001100" &
		"00001100" &
		"00000000" &
		"00000000" &

		"11000110" &
		"11001100" &
		"11011000" &
		"00111111" &
		"01100011" &
		"11001111" &
		"10001100" &
		"00001111" &

		"11000011" &
		"11000110" &
		"11001100" &
		"11011011" &
		"00110111" &
		"01101101" &
		"11001111" &
		"00000011" &

		"00011000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00000000" &
		"00110011" &
		"01100110" &
		"11001100" &
		"01100110" &
		"00110011" &
		"00000000" &
		"00000000" &

		"00000000" &
		"11001100" &
		"01100110" &
		"00110011" &
		"01100110" &
		"11001100" &
		"00000000" &
		"00000000" &

		"00100010" &
		"10001000" &
		"00100010" &
		"10001000" &
		"00100010" &
		"10001000" &
		"00100010" &
		"10001000" &

		"01010101" &
		"10101010" &
		"01010101" &
		"10101010" &
		"01010101" &
		"10101010" &
		"01010101" &
		"10101010" &

		"11011101" &
		"01110111" &
		"11011101" &
		"01110111" &
		"11011101" &
		"01110111" &
		"11011101" &
		"01110111" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"11111000" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00011000" &
		"00011000" &
		"11111000" &
		"00011000" &
		"11111000" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"11110110" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111110" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00000000" &
		"00000000" &
		"11111000" &
		"00011000" &
		"11111000" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00110110" &
		"00110110" &
		"11110110" &
		"00000110" &
		"11110110" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00000000" &
		"00000000" &
		"11111110" &
		"00000110" &
		"11110110" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00110110" &
		"00110110" &
		"11110110" &
		"00000110" &
		"11111110" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"11111110" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"11111000" &
		"00011000" &
		"11111000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111000" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"11111111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111111" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011111" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"11111111" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00011000" &
		"00011000" &
		"00011111" &
		"00011000" &
		"00011111" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"00110111" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00110110" &
		"00110110" &
		"00110111" &
		"00110000" &
		"00111111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00111111" &
		"00110000" &
		"00110111" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00110110" &
		"00110110" &
		"11110111" &
		"00000000" &
		"11111111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11111111" &
		"00000000" &
		"11110111" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00110110" &
		"00110110" &
		"00110111" &
		"00110000" &
		"00110111" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00000000" &
		"00000000" &
		"11111111" &
		"00000000" &
		"11111111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00110110" &
		"00110110" &
		"11110111" &
		"00000000" &
		"11110111" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00011000" &
		"00011000" &
		"11111111" &
		"00000000" &
		"11111111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"11111111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11111111" &
		"00000000" &
		"11111111" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111111" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"00111111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011111" &
		"00011000" &
		"00011111" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00011111" &
		"00011000" &
		"00011111" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00111111" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00110110" &
		"00110110" &
		"00110110" &
		"00110110" &
		"11111111" &
		"00110110" &
		"00110110" &
		"00110110" &

		"00011000" &
		"00011000" &
		"11111111" &
		"00011000" &
		"11111111" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"11111000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00011111" &
		"00011000" &
		"00011000" &
		"00011000" &

		"11111111" &
		"11111111" &
		"11111111" &
		"11111111" &
		"11111111" &
		"11111111" &
		"11111111" &
		"11111111" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111111" &
		"11111111" &
		"11111111" &
		"11111111" &

		"11110000" &
		"11110000" &
		"11110000" &
		"11110000" &
		"11110000" &
		"11110000" &
		"11110000" &
		"11110000" &

		"00001111" &
		"00001111" &
		"00001111" &
		"00001111" &
		"00001111" &
		"00001111" &
		"00001111" &
		"00001111" &

		"11111111" &
		"11111111" &
		"11111111" &
		"11111111" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01110110" &
		"11011100" &
		"11001000" &
		"11011100" &
		"01110110" &
		"00000000" &

		"00111000" &
		"01101100" &
		"01101100" &
		"01111000" &
		"01101100" &
		"01100110" &
		"01101100" &
		"01100000" &

		"00000000" &
		"11111110" &
		"11000110" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11111110" &
		"01101100" &
		"01101100" &
		"01101100" &
		"01101100" &
		"00000000" &

		"11111110" &
		"01100000" &
		"00110000" &
		"00011000" &
		"00110000" &
		"01100000" &
		"11111110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"11011000" &
		"11011000" &
		"11011000" &
		"01110000" &
		"00000000" &

		"00000000" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01111100" &
		"01100000" &
		"11000000" &

		"00000000" &
		"01110110" &
		"11011100" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"01111110" &
		"00011000" &
		"00111100" &
		"01100110" &
		"01100110" &
		"00111100" &
		"00011000" &
		"01111110" &

		"00111100" &
		"01100110" &
		"11000011" &
		"11111111" &
		"11000011" &
		"01100110" &
		"00111100" &
		"00000000" &

		"00111100" &
		"01100110" &
		"11000011" &
		"11000011" &
		"01100110" &
		"01100110" &
		"11100111" &
		"00000000" &

		"00001110" &
		"00011000" &
		"00001100" &
		"01111110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"11011011" &
		"11011011" &
		"01111110" &
		"00000000" &
		"00000000" &

		"00000110" &
		"00001100" &
		"01111110" &
		"11011011" &
		"11011011" &
		"01111110" &
		"01100000" &
		"11000000" &

		"00111000" &
		"01100000" &
		"11000000" &
		"11111000" &
		"11000000" &
		"01100000" &
		"00111000" &
		"00000000" &

		"01111000" &
		"11001100" &
		"11001100" &
		"11001100" &
		"11001100" &
		"11001100" &
		"11001100" &
		"00000000" &

		"00000000" &
		"01111110" &
		"00000000" &
		"01111110" &
		"00000000" &
		"01111110" &
		"00000000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"01111110" &
		"00011000" &
		"00011000" &
		"00000000" &
		"01111110" &
		"00000000" &

		"01100000" &
		"00110000" &
		"00011000" &
		"00110000" &
		"01100000" &
		"00000000" &
		"11111100" &
		"00000000" &

		"00011000" &
		"00110000" &
		"01100000" &
		"00110000" &
		"00011000" &
		"00000000" &
		"11111100" &
		"00000000" &

		"00001110" &
		"00011011" &
		"00011011" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"11011000" &
		"11011000" &
		"01110000" &

		"00011000" &
		"00011000" &
		"00000000" &
		"01111110" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00000000" &
		"01110110" &
		"11011100" &
		"00000000" &
		"01110110" &
		"11011100" &
		"00000000" &
		"00000000" &

		"00111000" &
		"01101100" &
		"01101100" &
		"00111000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00001111" &
		"00001100" &
		"00001100" &
		"00001100" &
		"11101100" &
		"01101100" &
		"00111100" &
		"00011100" &

		"01111000" &
		"01101100" &
		"01101100" &
		"01101100" &
		"01101100" &
		"00000000" &
		"00000000" &
		"00000000" &

		"01111100" &
		"00001100" &
		"01111100" &
		"01100000" &
		"01111100" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00111100" &
		"00111100" &
		"00111100" &
		"00111100" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00010000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000");

	constant psf1mag32x16 : std_logic_vector(0 to 32*32*16-1) := (
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0001111111100000" &
		"0011111111110000" &
		"0111110011111000" &
		"1111100001111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111100001111100" &
		"0111110011111000" &
		"0011111111110000" &
		"0001111111100000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000001111000000" &
		"0000011111000000" &
		"0000111111000000" &
		"0001111111000000" &
		"0011111111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0011111111111100" &
		"0011111111111100" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0011111111110000" &
		"0111111111111000" &
		"1111100001111100" &
		"1111000000111100" &
		"1110000000111100" &
		"0000000000111100" &
		"0000000001111100" &
		"0000000011111000" &
		"0000000111110000" &
		"0000001111100000" &
		"0000011111000000" &
		"0000111110000000" &
		"0001111100000000" &
		"0011111000000000" &
		"0111110000000000" &
		"1111100000000000" &
		"1111000000111100" &
		"1111000000111100" &
		"1111111111111100" &
		"1111111111111100" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0011111111110000" &
		"0111111111111000" &
		"1111100001111100" &
		"1111000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000001111000" &
		"0000111111110000" &
		"0000111111110000" &
		"0000000001111000" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"1111000000111100" &
		"1111100001111100" &
		"0111111111111000" &
		"0011111111110000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000011110000" &
		"0000000111110000" &
		"0000001111110000" &
		"0000011111110000" &
		"0000111111110000" &
		"0001111111110000" &
		"0011111011110000" &
		"0111110011110000" &
		"1111100011110000" &
		"1111000011110000" &
		"1111111111111100" &
		"1111111111111100" &
		"0000000011110000" &
		"0000000011110000" &
		"0000000011110000" &
		"0000000011110000" &
		"0000000011110000" &
		"0000000011110000" &
		"0000001111111100" &
		"0000001111111100" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"1111111111111100" &
		"1111111111111100" &
		"1111000000000000" &
		"1111000000000000" &
		"1111000000000000" &
		"1111000000000000" &
		"1111000000000000" &
		"1111000000000000" &
		"1111111111110000" &
		"1111111111111000" &
		"0000000001111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"1111000000111100" &
		"1111100001111100" &
		"0111111111111000" &
		"0011111111110000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000111111110000" &
		"0001111111110000" &
		"0011111000000000" &
		"0111110000000000" &
		"1111100000000000" &
		"1111000000000000" &
		"1111000000000000" &
		"1111000000000000" &
		"1111111111110000" &
		"1111111111111000" &
		"1111100001111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111100001111100" &
		"0111111111111000" &
		"0011111111110000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"1111111111111100" &
		"1111111111111100" &
		"1111000000111100" &
		"1111000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000001111100" &
		"0000000011111000" &
		"0000000111110000" &
		"0000001111100000" &
		"0000011111000000" &
		"0000111110000000" &
		"0000111100000000" &
		"0000111100000000" &
		"0000111100000000" &
		"0000111100000000" &
		"0000111100000000" &
		"0000111100000000" &
		"0000111100000000" &
		"0000111100000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0011111111110000" &
		"0111111111111000" &
		"1111100001111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"0111100001111000" &
		"0011111111110000" &
		"0011111111110000" &
		"0111100001111000" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111100001111100" &
		"0111111111111000" &
		"0011111111110000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0011111111110000" &
		"0111111111111000" &
		"1111100001111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111100001111100" &
		"0111111111111100" &
		"0011111111111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000000111100" &
		"0000000001111100" &
		"0000000011111000" &
		"0000000111110000" &
		"0011111111100000" &
		"0011111111000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000001111000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000011110000000" &
		"0000011110000000" &
		"0000011110000000" &
		"0000011110000000" &
		"0111111111111000" &
		"0111111111111000" &
		"0111111111111000" &
		"0000011110000000" &
		"0000011110000000" &
		"0000011110000000" &
		"0000011110000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"1111111111111100" &
		"1111111111111100" &
		"1111111111111100" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"1111110011110000" &
		"1111111111111000" &
		"1111111111111100" &
		"1111111111111100" &
		"1111001100111100" &
		"1111001100111100" &
		"1111001100111100" &
		"1111001100111100" &
		"1111001100111100" &
		"1111001100111100" &
		"1111001100111100" &
		"1111001100111100" &
		"1111000000111100" &
		"1111000000111100" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &


		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011111111111000" &
		"0011111111110000" &
		"0011110000000000" &
		"0011110000000000" &
		"0011110000000000" &
		"0011110000000000" &
		"1111100000000000" &
		"1111000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"1111001111110000" &
		"1111111111111000" &
		"0011111001111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0011110000111100" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0011111111110000" &
		"0111111111111000" &
		"1111000001111100" &
		"1111000000111100" &
		"0111100000000000" &
		"0011111000000000" &
		"0001111110000000" &
		"0000011111100000" &
		"0000000111110000" &
		"0000000001111000" &
		"1111000000111100" &
		"1111100000111100" &
		"0111111111111000" &
		"0011111111110000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111000000111100" &
		"1111100001111100" &
		"0111110011111000" &
		"0011111111110000" &
		"0001111111100000" &
		"0000111111000000" &
		"0000011110000000" &
		"0000001100000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &
		"0000000000000000" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------");

	constant psf1hex8x16 : std_logic_vector(0 to 16*8*16-1) := (
		-- x"30" --
		"00000000" & --"00000000" &
		"00000000" & --"00000000" &
		"00000000" & --"00111000" &
		"00000000" & --"01101100" &
		"00000000" & --"11000110" &
		"00000000" & --"11000110" &
		"00000000" & --"11010110" &
		"00000000" & --"11010110" &
		"00000000" & --"11000110" &
		"00000000" & --"11000110" &
		"00000000" & --"01101100" &
		"00000000" & --"00111000" &
		"00000000" & --"00000000" &
		"00000000" & --"00000000" &
		"00000000" & --"00000000" &
		"00000000" & --"00000000" &

		-- x"31" --
		"00000000" &
		"00000000" &
		"00011000" &
		"00111000" &
		"01111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"32" --
		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"01100000" &
		"11000000" &
		"11000110" &
		"11111110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"33" --
		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"00000110" &
		"00000110" &
		"00111100" &
		"00000110" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"34" --
		"00000000" &
		"00000000" &
		"00001100" &
		"00011100" &
		"00111100" &
		"01101100" &
		"11001100" &
		"11111110" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00011110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"35" --
		"00000000" &
		"00000000" &
		"11111110" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11111100" &
		"00000110" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"36" --
		"00000000" &
		"00000000" &
		"00111000" &
		"01100000" &
		"11000000" &
		"11000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"37" --
		"00000000" &
		"00000000" &
		"11111110" &
		"11000110" &
		"00000110" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"38" --
		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"39" --
		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"00000110" &
		"00000110" &
		"00001100" &
		"01111000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"41" --
		"00000000" &
		"00000000" &
		"00010000" &
		"00111000" &
		"01101100" &
		"11000110" &
		"11000110" &
		"11111110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"42" --
		"00000000" &
		"00000000" &
		"11111100" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01111100" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"11111100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"43" --
		"00000000" &
		"00000000" &
		"00111100" &
		"01100110" &
		"11000010" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000010" &
		"01100110" &
		"00111100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"44" --
		"00000000" &
		"00000000" &
		"11111000" &
		"01101100" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01101100" &
		"11111000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"45" --
		"00000000" &
		"00000000" &
		"11111110" &
		"01100110" &
		"01100010" &
		"01101000" &
		"01111000" &
		"01101000" &
		"01100000" &
		"01100010" &
		"01100110" &
		"11111110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		-- x"46" --
		"00000000" &
		"00000000" &
		"11111110" &
		"01100110" &
		"01100010" &
		"01101000" &
		"01111000" &
		"01101000" &
		"01100000" &
		"01100000" &
		"01100000" &
		"11110000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000");

	function shuffle_code (
		constant font   : std_logic_vector;
		constant width  : natural;
		constant height : natural)
		return std_logic_vector;
end;

package body cgafonts is

	function shuffle_code (
		constant font   : std_logic_vector;
		constant width  : natural;
		constant height : natural)
		return std_logic_vector is
		variable retval : std_logic_vector(font'range) := (others => '-');
		constant codes  : natural := font'length/(width*height);
	begin
		for k in 0 to codes-1 loop
			for i in 0 to height-1 loop
				for j in 0 to width-1 loop
					retval(codes*(width*i+j)+k) := font(width*(height*k+i)+j);
				end loop;
			end loop;
		end loop;
		return retval;
	end;
end;

