library foo;
use foo.test.all;

entity due is
end;

architecture def of due is
begin
	process
		variable myvar : natural;
		variable mesg  : std.textio.line;
	begin
		myvar := std;
	end process;
end;
