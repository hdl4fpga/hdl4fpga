library ieee;
use ieee.std_logic_1164.all;

package cgafonts3 is

                                    
constant psf1cp850x8x16_00_to_F7 : std_logic_vector(0 to 128*8*16-1) := (

		-- xB"00" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"01" --
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"10000001" &
		B"10100101" &
		B"10000001" &
		B"10000001" &
		B"10111101" &
		B"10011001" &
		B"10000001" &
		B"10000001" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"02" --
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"11111111" &
		B"11011011" &
		B"11111111" &
		B"11111111" &
		B"11000011" &
		B"11100111" &
		B"11111111" &
		B"11111111" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"03" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01101100" &
		B"11111110" &
		B"11111110" &
		B"11111110" &
		B"11111110" &
		B"01111100" &
		B"00111000" &
		B"00010000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"04" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01111100" &
		B"11111110" &
		B"01111100" &
		B"00111000" &
		B"00010000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"05" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"00111100" &
		B"11100111" &
		B"11100111" &
		B"11100111" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"06" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"11111111" &
		B"11111111" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"07" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"00111100" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"08" --
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11100111" &
		B"11000011" &
		B"11000011" &
		B"11100111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &

		-- xB"09" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"01100110" &
		B"01000010" &
		B"01000010" &
		B"01100110" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"0a" --
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11000011" &
		B"10011001" &
		B"10111101" &
		B"10111101" &
		B"10011001" &
		B"11000011" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &

		-- xB"0b" --
		B"00000000" &
		B"00000000" &
		B"00011110" &
		B"00001110" &
		B"00011010" &
		B"00110010" &
		B"01111000" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"0c" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"0d" --
		B"00000000" &
		B"00000000" &
		B"00111111" &
		B"00110011" &
		B"00111111" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"01110000" &
		B"11110000" &
		B"11100000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"0e" --
		B"00000000" &
		B"00000000" &
		B"01111111" &
		B"01100011" &
		B"01111111" &
		B"01100011" &
		B"01100011" &
		B"01100011" &
		B"01100011" &
		B"01100111" &
		B"11100111" &
		B"11100110" &
		B"11000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"0f" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"11011011" &
		B"00111100" &
		B"11100111" &
		B"00111100" &
		B"11011011" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"10" --
		B"00000000" &
		B"10000000" &
		B"11000000" &
		B"11100000" &
		B"11110000" &
		B"11111000" &
		B"11111110" &
		B"11111000" &
		B"11110000" &
		B"11100000" &
		B"11000000" &
		B"10000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"11" --
		B"00000000" &
		B"00000010" &
		B"00000110" &
		B"00001110" &
		B"00011110" &
		B"00111110" &
		B"11111110" &
		B"00111110" &
		B"00011110" &
		B"00001110" &
		B"00000110" &
		B"00000010" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"12" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00111100" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"13" --
		B"00000000" &
		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"14" --
		B"00000000" &
		B"00000000" &
		B"01111111" &
		B"11011011" &
		B"11011011" &
		B"11011011" &
		B"01111011" &
		B"00011011" &
		B"00011011" &
		B"00011011" &
		B"00011011" &
		B"00011011" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"15" --
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"01100000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"00001100" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"16" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"11111110" &
		B"11111110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"17" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00111100" &
		B"00011000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"18" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"19" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00111100" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"1a" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00001100" &
		B"11111110" &
		B"00001100" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"1b" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00110000" &
		B"01100000" &
		B"11111110" &
		B"01100000" &
		B"00110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"1c" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"1d" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00101000" &
		B"01101100" &
		B"11111110" &
		B"01101100" &
		B"00101000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"1e" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"00111000" &
		B"01111100" &
		B"01111100" &
		B"11111110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- xB"1f" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"11111110" &
		B"01111100" &
		B"01111100" &
		B"00111000" &
		B"00111000" &
		B"00010000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"20" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"21" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"00111100" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"22" --
		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00100100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"23" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01101100" &
		B"01101100" &
		B"11111110" &
		B"01101100" &
		B"01101100" &
		B"01101100" &
		B"11111110" &
		B"01101100" &
		B"01101100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"24" --
		B"00011000" &
		B"00011000" &
		B"01111100" &
		B"11000110" &
		B"11000010" &
		B"11000000" &
		B"01111100" &
		B"00000110" &
		B"00000110" &
		B"10000110" &
		B"11000110" &
		B"01111100" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &

		-- x"25" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11000010" &
		B"11000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11000110" &
		B"10000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"26" --
		B"00000000" &
		B"00000000" &
		B"00111000" &
		B"01101100" &
		B"01101100" &
		B"00111000" &
		B"01110110" &
		B"11011100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"27" --
		B"00000000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"01100000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"28" --
		B"00000000" &
		B"00000000" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"29" --
		B"00000000" &
		B"00000000" &
		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"2a" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01100110" &
		B"00111100" &
		B"11111111" &
		B"00111100" &
		B"01100110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"2b" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"2c" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"2d" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"2e" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"2f" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000010" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11000000" &
		B"10000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"30" --
		B"00000000" &
		B"00000000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11010110" &
		B"11010110" &
		B"11000110" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"31" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111000" &
		B"01111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"32" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11000000" &
		B"11000110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"33" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"00000110" &
		B"00000110" &
		B"00111100" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"34" --
		B"00000000" &
		B"00000000" &
		B"00001100" &
		B"00011100" &
		B"00111100" &
		B"01101100" &
		B"11001100" &
		B"11111110" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00011110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"35" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11111100" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"36" --
		B"00000000" &
		B"00000000" &
		B"00111000" &
		B"01100000" &
		B"11000000" &
		B"11000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"37" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"11000110" &
		B"00000110" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"38" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"39" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00001100" &
		B"01111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"3a" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"3b" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"3c" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"3d" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"3e" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"3f" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"00001100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"40" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11011110" &
		B"11011110" &
		B"11011110" &
		B"11011100" &
		B"11000000" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"41" --
		B"00000000" &
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"42" --
		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"11111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"43" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"01100110" &
		B"11000010" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000010" &
		B"01100110" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"44" --
		B"00000000" &
		B"00000000" &
		B"11111000" &
		B"01101100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01101100" &
		B"11111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"45" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"01100110" &
		B"01100010" &
		B"01101000" &
		B"01111000" &
		B"01101000" &
		B"01100000" &
		B"01100010" &
		B"01100110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"46" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"01100110" &
		B"01100010" &
		B"01101000" &
		B"01111000" &
		B"01101000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"11110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"47" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"01100110" &
		B"11000010" &
		B"11000000" &
		B"11000000" &
		B"11011110" &
		B"11000110" &
		B"11000110" &
		B"01100110" &
		B"00111010" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"48" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"49" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"4a" --
		B"00000000" &
		B"00000000" &
		B"00011110" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"4b" --
		B"00000000" &
		B"00000000" &
		B"11100110" &
		B"01100110" &
		B"01100110" &
		B"01101100" &
		B"01111000" &
		B"01111000" &
		B"01101100" &
		B"01100110" &
		B"01100110" &
		B"11100110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"4c" --
		B"00000000" &
		B"00000000" &
		B"11110000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"01100010" &
		B"01100110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"4d" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11101110" &
		B"11111110" &
		B"11111110" &
		B"11010110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"4e" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11100110" &
		B"11110110" &
		B"11111110" &
		B"11011110" &
		B"11001110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"4f" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"50" --
		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"11110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"51" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11010110" &
		B"11011110" &
		B"01111100" &
		B"00001100" &
		B"00001110" &
		B"00000000" &
		B"00000000" &

		-- x"52" --
		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01101100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"11100110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"53" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"01100000" &
		B"00111000" &
		B"00001100" &
		B"00000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"54" --
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"01111110" &
		B"01011010" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"55" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"56" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"00010000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"57" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11010110" &
		B"11010110" &
		B"11010110" &
		B"11111110" &
		B"11101110" &
		B"01101100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"58" --
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"01101100" &
		B"01111100" &
		B"00111000" &
		B"00111000" &
		B"01111100" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"59" --
		B"00000000" &
		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"5a" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"11000110" &
		B"10000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11000010" &
		B"11000110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"5b" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"5c" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"10000000" &
		B"11000000" &
		B"11100000" &
		B"01110000" &
		B"00111000" &
		B"00011100" &
		B"00001110" &
		B"00000110" &
		B"00000010" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"5d" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"5e" --
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"5f" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &

		-- x"60" --
		B"00000000" &
		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"61" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111000" &
		B"00001100" &
		B"01111100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"62" --
		B"00000000" &
		B"00000000" &
		B"11100000" &
		B"01100000" &
		B"01100000" &
		B"01111000" &
		B"01101100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"63" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"64" --
		B"00000000" &
		B"00000000" &
		B"00011100" &
		B"00001100" &
		B"00001100" &
		B"00111100" &
		B"01101100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"65" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"66" --
		B"00000000" &
		B"00000000" &
		B"00011100" &
		B"00110110" &
		B"00110010" &
		B"00110000" &
		B"01111000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"01111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"67" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01110110" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01111100" &
		B"00001100" &
		B"11001100" &
		B"01111000" &
		B"00000000" &

		-- x"68" --
		B"00000000" &
		B"00000000" &
		B"11100000" &
		B"01100000" &
		B"01100000" &
		B"01101100" &
		B"01110110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"11100110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"69" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"6a" --
		B"00000000" &
		B"00000000" &
		B"00000110" &
		B"00000110" &
		B"00000000" &
		B"00001110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00000000" &

		-- x"6b" --
		B"00000000" &
		B"00000000" &
		B"11100000" &
		B"01100000" &
		B"01100000" &
		B"01100110" &
		B"01101100" &
		B"01111000" &
		B"01111000" &
		B"01101100" &
		B"01100110" &
		B"11100110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"6c" --
		B"00000000" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"6d" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11101100" &
		B"11111110" &
		B"11010110" &
		B"11010110" &
		B"11010110" &
		B"11010110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"6e" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11011100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"6f" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"70" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11011100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01100000" &
		B"01100000" &
		B"11110000" &
		B"00000000" &

		-- x"71" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01110110" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01111100" &
		B"00001100" &
		B"00001100" &
		B"00011110" &
		B"00000000" &

		-- x"72" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11011100" &
		B"01110110" &
		B"01100110" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"11110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"73" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"01100000" &
		B"00111000" &
		B"00001100" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"74" --
		B"00000000" &
		B"00000000" &
		B"00010000" &
		B"00110000" &
		B"00110000" &
		B"11111100" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110110" &
		B"00011100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"75" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"76" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"77" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11010110" &
		B"11010110" &
		B"11010110" &
		B"11111110" &
		B"01101100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"78" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"00111000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"79" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"00001100" &
		B"11111000" &
		B"00000000" &

		-- x"7a" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"11001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11000110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"7b" --
		B"00000000" &
		B"00000000" &
		B"00001110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01110000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00001110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"7c" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"7d" --
		B"00000000" &
		B"00000000" &
		B"01110000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00001110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"7e" --
		B"00000000" &
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"7f" --
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000"
		);

end;
