-- (c) EMARD
-- License=BSD

library ieee;
use ieee.std_logic_1164.all;

-- OLED FONT

package oled_font_pack is
  type T_oled_char is array (0 to 7) of std_logic_vector(4 downto 0);
  type T_oled_font is array (0 to 16) of T_oled_char;
  constant C_oled_font: T_oled_font :=
  (
    ( -- 0
      "01110",
      "10001",
      "10011",
      "10101",
      "11001",
      "10001",
      "01110",
      "00000"
    ),
    ( -- 1
      "00100",
      "01100",
      "00100",
      "00100",
      "00100",
      "00100",
      "01110",
      "00000"
    ),
    ( -- 2
      "01110",
      "10001",
      "00001",
      "00010",
      "00100",
      "01000",
      "11111",
      "00000"
    ),
    ( -- 3
      "01110",
      "10001",
      "00001",
      "01110",
      "00001",
      "10001",
      "01110",
      "00000"
    ),
    ( -- 4
      "00010",
      "00110",
      "01010",
      "10010",
      "11111",
      "00010",
      "00010",
      "00000"
    ),
    ( -- 5
      "11111",
      "10000",
      "11110",
      "00001",
      "00001",
      "10001",
      "01110",
      "00000"
    ),
    ( -- 6
      "01111",
      "10000",
      "11110",
      "10001",
      "10001",
      "10001",
      "01110",
      "00000"
    ),
    ( -- 7
      "11111",
      "10001",
      "00001",
      "00010",
      "00100",
      "01000",
      "01000",
      "00000"
    ),
    ( -- 8
      "01110",
      "10001",
      "10001",
      "01110",
      "10001",
      "10001",
      "01110",
      "00000"
    ),
    ( -- 9
      "01110",
      "10001",
      "10001",
      "01111",
      "00001",
      "10001",
      "01110",
      "00000"
    ),
    ( -- 10: A
      "01110",
      "10001",
      "10001",
      "11111",
      "10001",
      "10001",
      "10001",
      "00000"
    ),
    ( -- 11: B
      "11110",
      "10001",
      "10001",
      "11110",
      "10001",
      "10001",
      "11110",
      "00000"
    ),
    ( -- 12: C
      "01110",
      "10001",
      "10000",
      "10000",
      "10000",
      "10001",
      "01110",
      "00000"
    ),
    ( -- 13: D
      "11110",
      "10001",
      "10001",
      "10001",
      "10001",
      "10001",
      "11110",
      "00000"
    ),
    ( -- 14: E
      "11111",
      "10000",
      "10000",
      "11110",
      "10000",
      "10000",
      "11111",
      "00000"
    ),
    ( -- 15: F
      "11111",
      "10000",
      "10000",
      "11110",
      "10000",
      "10000",
      "10000",
      "00000"
    ),
    ( -- 16: SPACE
      "00000",
      "00000",
      "00000",
      "00000",
      "00000",
      "00000",
      "00000",
      "00000"
    )
  );
end;
