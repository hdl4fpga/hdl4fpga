--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library hdl4fpga;
use  hdl4fpga.std.all;
use  hdl4fpga.scopeiopkg.all;

architecture scopeiopkg of testbench is

		constant width  : natural := 33;
		constant height : natural := 10;
		constant layout : tag_vector(analogtime_layout'range) := text_setaddr(
			analogtime_layout, 
			width,
			height);
		constant rom    : std_logic_vector(0 to width*height*ascii'length-1) := text_content(
			analogtime_layout, 
			width,
			height,
			lang_en);
begin

	process
		variable mesg : line;
	begin
		wait;
	end process;

end;
