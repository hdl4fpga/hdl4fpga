library ieee;
use ieee.std_logic_1164.all;

package cgafonts7 is

	constant psf1mag32x16 : std_logic_vector(0 to 32*32*16-1) := (
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0001111111100000" &
		B"0011111111110000" &
		B"0111110011111000" &
		B"1111100001111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111100001111100" &
		B"0111110011111000" &
		B"0011111111110000" &
		B"0001111111100000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000001111000000" &
		B"0000011111000000" &
		B"0000111111000000" &
		B"0001111111000000" &
		B"0011111111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0011111111111100" &
		B"0011111111111100" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0011111111110000" &
		B"0111111111111000" &
		B"1111100001111100" &
		B"1111000000111100" &
		B"1110000000111100" &
		B"0000000000111100" &
		B"0000000001111100" &
		B"0000000011111000" &
		B"0000000111110000" &
		B"0000001111100000" &
		B"0000011111000000" &
		B"0000111110000000" &
		B"0001111100000000" &
		B"0011111000000000" &
		B"0111110000000000" &
		B"1111100000000000" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111111111111100" &
		B"1111111111111100" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0011111111110000" &
		B"0111111111111000" &
		B"1111100001111100" &
		B"1111000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000001111000" &
		B"0000111111110000" &
		B"0000111111110000" &
		B"0000000001111000" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"1111000000111100" &
		B"1111100001111100" &
		B"0111111111111000" &
		B"0011111111110000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000011110000" &
		B"0000000111110000" &
		B"0000001111110000" &
		B"0000011111110000" &
		B"0000111111110000" &
		B"0001111111110000" &
		B"0011111011110000" &
		B"0111110011110000" &
		B"1111100011110000" &
		B"1111000011110000" &
		B"1111111111111100" &
		B"1111111111111100" &
		B"0000000011110000" &
		B"0000000011110000" &
		B"0000000011110000" &
		B"0000000011110000" &
		B"0000000011110000" &
		B"0000000011110000" &
		B"0000001111111100" &
		B"0000001111111100" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"1111111111111100" &
		B"1111111111111100" &
		B"1111000000000000" &
		B"1111000000000000" &
		B"1111000000000000" &
		B"1111000000000000" &
		B"1111000000000000" &
		B"1111000000000000" &
		B"1111111111110000" &
		B"1111111111111000" &
		B"0000000001111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"1111000000111100" &
		B"1111100001111100" &
		B"0111111111111000" &
		B"0011111111110000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000111111110000" &
		B"0001111111110000" &
		B"0011111000000000" &
		B"0111110000000000" &
		B"1111100000000000" &
		B"1111000000000000" &
		B"1111000000000000" &
		B"1111000000000000" &
		B"1111111111110000" &
		B"1111111111111000" &
		B"1111100001111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111100001111100" &
		B"0111111111111000" &
		B"0011111111110000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"1111111111111100" &
		B"1111111111111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000001111100" &
		B"0000000011111000" &
		B"0000000111110000" &
		B"0000001111100000" &
		B"0000011111000000" &
		B"0000111110000000" &
		B"0000111100000000" &
		B"0000111100000000" &
		B"0000111100000000" &
		B"0000111100000000" &
		B"0000111100000000" &
		B"0000111100000000" &
		B"0000111100000000" &
		B"0000111100000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0011111111110000" &
		B"0111111111111000" &
		B"1111100001111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"0111100001111000" &
		B"0011111111110000" &
		B"0011111111110000" &
		B"0111100001111000" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111100001111100" &
		B"0111111111111000" &
		B"0011111111110000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0011111111110000" &
		B"0111111111111000" &
		B"1111100001111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111100001111100" &
		B"0111111111111100" &
		B"0011111111111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000000111100" &
		B"0000000001111100" &
		B"0000000011111000" &
		B"0000000111110000" &
		B"0011111111100000" &
		B"0011111111000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000001111000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000011110000000" &
		B"0000011110000000" &
		B"0000011110000000" &
		B"0000011110000000" &
		B"0111111111111000" &
		B"0111111111111000" &
		B"0111111111111000" &
		B"0000011110000000" &
		B"0000011110000000" &
		B"0000011110000000" &
		B"0000011110000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"1111111111111100" &
		B"1111111111111100" &
		B"1111111111111100" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"1111110011110000" &
		B"1111111111111000" &
		B"1111111111111100" &
		B"1111111111111100" &
		B"1111001100111100" &
		B"1111001100111100" &
		B"1111001100111100" &
		B"1111001100111100" &
		B"1111001100111100" &
		B"1111001100111100" &
		B"1111001100111100" &
		B"1111001100111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &


		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011111111111000" &
		B"0011111111110000" &
		B"0011110000000000" &
		B"0011110000000000" &
		B"0011110000000000" &
		B"0011110000000000" &
		B"1111100000000000" &
		B"1111000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"1111001111110000" &
		B"1111111111111000" &
		B"0011111001111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0011110000111100" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0011111111110000" &
		B"0111111111111000" &
		B"1111000001111100" &
		B"1111000000111100" &
		B"0111100000000000" &
		B"0011111000000000" &
		B"0001111110000000" &
		B"0000011111100000" &
		B"0000000111110000" &
		B"0000000001111000" &
		B"1111000000111100" &
		B"1111100000111100" &
		B"0111111111111000" &
		B"0011111111110000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111000000111100" &
		B"1111100001111100" &
		B"0111110011111000" &
		B"0011111111110000" &
		B"0001111111100000" &
		B"0000111111000000" &
		B"0000011110000000" &
		B"0000001100000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &
		B"0000000000000000" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &

		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------" &
		"----------------");

	constant psf1hex8x16 : std_logic_vector(0 to 16*8*16-1) := (
		-- x"30" --
		B"00000000" & --B"00000000" &
		B"00000000" & --B"00000000" &
		B"00000000" & --B"00111000" &
		B"00000000" & --B"01101100" &
		B"00000000" & --B"11000110" &
		B"00000000" & --B"11000110" &
		B"00000000" & --B"11010110" &
		B"00000000" & --B"11010110" &
		B"00000000" & --B"11000110" &
		B"00000000" & --B"11000110" &
		B"00000000" & --B"01101100" &
		B"00000000" & --B"00111000" &
		B"00000000" & --B"00000000" &
		B"00000000" & --B"00000000" &
		B"00000000" & --B"00000000" &
		B"00000000" & --B"00000000" &

		-- x"31" --
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111000" &
		B"01111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"32" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11000000" &
		B"11000110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"33" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"00000110" &
		B"00000110" &
		B"00111100" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"34" --
		B"00000000" &
		B"00000000" &
		B"00001100" &
		B"00011100" &
		B"00111100" &
		B"01101100" &
		B"11001100" &
		B"11111110" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00011110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"35" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11111100" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"36" --
		B"00000000" &
		B"00000000" &
		B"00111000" &
		B"01100000" &
		B"11000000" &
		B"11000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"37" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"11000110" &
		B"00000110" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"38" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"39" --
		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00001100" &
		B"01111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"41" --
		B"00000000" &
		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"42" --
		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"11111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"43" --
		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"01100110" &
		B"11000010" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000010" &
		B"01100110" &
		B"00111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"44" --
		B"00000000" &
		B"00000000" &
		B"11111000" &
		B"01101100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01101100" &
		B"11111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"45" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"01100110" &
		B"01100010" &
		B"01101000" &
		B"01111000" &
		B"01101000" &
		B"01100000" &
		B"01100010" &
		B"01100110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		-- x"46" --
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"01100110" &
		B"01100010" &
		B"01101000" &
		B"01111000" &
		B"01101000" &
		B"01100000" &
		B"01100000" &
		B"01100000" &
		B"11110000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000");

end;
