use std.textio.all;

library foo;
use foo.test.all;

entity due is
	port (
		i : in std);
end;

