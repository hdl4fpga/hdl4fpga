library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity adjdll is
	port (
		rst  : in  std_logic;
		sclk : in  std_logic;
		eclk : in  std_logic;
		kclk : in  std_logic;
		stop : out std_logic;
		rdy  : out std_logic;
		pha  : out std_logic_vector);
		
end;

architecture beh of adjdll is

	signal ph : std_logic_vector(pha'range);
	signal qk : std_logic;
	signal ok : std_logic;
	signal prdy : std_logic_vector(0 to 4);

begin

	process (rst, kclk)
	begin
		if rst='1' then
			qk <= '0';
		elsif rising_edge(kclk) then
			qk <= not qk;
		end if;
	end process;

	process (rst, sclk)
		variable q : std_logic_vector(0 to 1);
	begin
		if rst='1' then
			ok <= '0';
			q := (others => '0');
		elsif rising_edge(sclk) then
			if prdy(0)='0' then
				ok <= not q(0) and q(1);
			end if;

			q(0) := eclk;
			q(1) := qk;
		end if;
	end process;

	process(rst, sclk)
		variable dg : unsigned(0 to pha'length+1);
		variable dy : unsigned(prdy'range);
		variable aux : unsigned(pha'range);
	begin
		if rst='1' then
			ph <= (others => '0');
			dg := (0 => '1', others => '0');
			rdy <= dg(dg'right);
			dy := (others => '0');
			prdy <= (others => '0');
		elsif rising_edge(sclk) then
			if dg(dg'right)='0' then
				if prdy(3)='1' then
					aux := unsigned(ph);
					aux := aux or dg(0 to ph'length-1);
					if ok='0' then
						aux := aux and not dg(1 to ph'length);
					end if;
					ph <= std_logic_vector(aux);
					dg := dg srl 1;
				end if;
				prdy <= std_logic_vector(dy and not (dy ror 1));
				dy := dy(1 to dy'right) & not dy(0);
			else
				prdy <= (others => '0');
			end if;
			rdy <= dg(dg'right);
		end if;
	end process;
	stop <= prdy(2);
	pha <= ph;
end;
