--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library hdl4fpga;
use hdl4fpga.std.all;

entity scopeio_axisticks is
	port (
		clk         : in  std_logic;

		axis_req    : in  std_logic;
		axis_rdy    : out std_logic;
		axis_unit   : in  std_logic_vector;
		axis_escale : in  std_logic_vector;

		hz_length   : in  std_logic_vector := b"110";
		hz_offset   : in  std_logic_vector;
		hz_dv       : out std_logic;

		vt_length   : in  std_logic_vector := b"100";
		vt_offset   : in  std_logic_vector := std_logic_vector'(b"0000");
		vt_dv       : out std_logic;

		tick        : out std_logic_vector;
		value       : out std_logic_vector);
end;

architecture def of scopeio_axisticks is

	signal wrt_req : std_logic;
	signal wrt_rdy : std_logic;
	signal wrt_length : std_logic_vector(0 to 3-1);

	signal bin_dv  : std_logic;
	signal bin_val : std_logic_vector(4*4-1 downto 0);
	signal bcd_dv  : std_logic;

	signal vt_gnt  : std_logic;
	signal hz_gnt  : std_logic;

	signal dev_req : std_logic_vector(1 to 2);
	signal dev_rdy : std_logic_vector(1 to 2);
	signal dev_gnt : std_logic_vector(1 to 2);

	signal base    : std_logic_vector(8-1 downto 0);
	signal from    : signed(base'range);
	signal unit    : unsigned(base'range);

begin

	from <= resize(  signed(axis_from), base'length);
	unit <= resize(unsigned(axis_unit), base'length);

	mult_b : block
		signal ini : std_logic; 
	begin
		ini <= '1';
		mult_e : entity hdl4fpga.mult
		port map (
			clk     => clk,
			ini     => ini,
			multand => std_logic_vector(from(4-1 downto 0)),
			multier => std_logic_vector(unit(4-1 downto 0)),
			product => base);
	end block;

	process(clk)
		variable cntr : signed(bin_val'range);
	begin
		if rising_edge(clk) then
			if wrt_req='0' then
				cntr := (others => '0');
			elsif wrt_rdy='0' then
				if bin_dv='1' then
					cntr := cntr + signed(axis_unit);
				end if;
			end if;
			if hz_gnt='1' then
				bin_val <= std_logic_vector((cntr + signed(base)) sll 1);
			else
				bin_val <= std_logic_vector(cntr + signed(base));
			end if;
		end if;
	end process;

	wrt_length <= wirebus(hz_length & vt_length, dev_gnt);

	scopeio_write_e : entity hdl4fpga.scopeio_writeticks
	port map (
		clk        => clk,
		write_req  => axis_req,
		write_rdy  => axis_rdy,
		point      => axis_point,
		length     => wrt_length,
		element    => tick,
		bin_dv     => bin_dv,
		bin_val    => bin_val,
		bcd_sign   => vt_gnt,
		bcd_left   => hz_gnt,
		bcd_dv     => bcd_dv,
		bcd_val    => value);

	hz_dv <= bcd_dv and hz_gnt;
	vt_dv <= bcd_dv and vt_gnt;

end;
