--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity xc7a_ddrdqphy is
	generic (
		taps      : natural;
		data_gear : natural;
		data_edge : boolean;
		byte_size : natural);
	port (
		tp_sel    : in  std_logic;
		tp_delay  : out std_logic_vector(8-1 downto 0);

		sys_rsts  : in  std_logic_vector;
		sys_clks  : in  std_logic_vector;
		sys_wlreq : in  std_logic;
		sys_wlrdy : out std_logic;
		sys_rlreq : in  std_logic;
		sys_rlrdy : buffer std_logic;
		sys_rlcal : out std_logic;
		sys_dmt   : in  std_logic_vector(0 to DATA_GEAR-1) := (others => '-');
		sys_dmi   : in  std_logic_vector(DATA_GEAR-1 downto 0) := (others => '-');
		sys_sti   : in  std_logic_vector(0 to DATA_GEAR-1) := (others => '-');
		sys_sto   : out std_logic_vector(0 to DATA_GEAR-1);
		sys_dqi   : in  std_logic_vector(DATA_GEAR*BYTE_SIZE-1 downto 0);
		sys_dqt   : in  std_logic_vector(DATA_GEAR-1 downto 0);
		sys_dqo   : out std_logic_vector(DATA_GEAR*BYTE_SIZE-1 downto 0);
		sys_dqso  : in  std_logic_vector(0 to DATA_GEAR-1);
		sys_dqst  : in  std_logic_vector(0 to DATA_GEAR-1);

		ddr_dmt   : out std_logic;
		ddr_dmo   : out std_logic;
		ddr_dqsi  : in  std_logic;
		ddr_dqi   : in  std_logic_vector(BYTE_SIZE-1 downto 0);
		ddr_dqt   : out std_logic_vector(BYTE_SIZE-1 downto 0);
		ddr_dqo   : out std_logic_vector(BYTE_SIZE-1 downto 0);

		ddr_dqst  : out std_logic;
		ddr_dqso  : out std_logic);

		constant clk0div  : natural := 0;
		constant clk90div : natural := 1;
		constant iodclk   : natural := 2;
		constant clk0     : natural := 3;
		constant clk90    : natural := 4;

		constant rst0div  : natural := 0;
		constant rst90div : natural := 1;
		constant rstiod   : natural := 1;
end;

library hdl4fpga;
use hdl4fpga.std.all;

architecture virtex7 of xc7a_ddrdqphy is

	signal adjdqs_req : std_logic;
	signal adjdqs_rdy : std_logic;
	signal adjdqi_req : std_logic;
	signal adjdqi_rdy : std_logic_vector(ddr_dqi'range);
	signal adjsto_req : std_logic;
	signal adjsto_rdy : std_logic;

	signal iod_rst    : std_logic;
	signal dqsi_buf   : std_logic;
	signal dqsiod_inc : std_logic;
	signal dqsiod_ce  : std_logic;

	signal dqs180     : std_logic;
	signal dqspre     : std_logic;
	signal dq         : std_logic_vector(sys_dqo'range);
	signal dqi        : std_logic_vector(ddr_dqi'range);
	signal dqh        : std_logic_vector(dq'range);
	signal dqf        : std_logic_vector(dq'range);

	signal tp_dqidly  : std_logic_vector(0 to 5-1);
	signal tp_dqsdly  : std_logic_vector(0 to 5-1);
	signal tp_dqssel  : std_logic_vector(0 to 3-1);

	constant dqs_linedelay : time := 1.35 ns;
	constant dqi_linedelay : time := 0 ns; --1.35 ns;

begin

	with tp_sel select
	tp_delay <=
		dqs180 & dqspre & std_logic_vector(resize(unsigned(tp_dqidly), tp_delay'length-2)) when '1',
		std_logic_vector(resize(unsigned(std_logic_vector'(tp_dqssel & tp_dqsdly)), tp_delay'length)) when others;

	sys_wlrdy <= sys_wlreq;

	process (sys_clks(iodclk))
		type states is (sync_start, sync_dqs, sync_dqi, sync_sto);
		variable state : states;
		variable aux : bit;
	begin
		if rising_edge(sys_clks(iodclk)) then
			if (to_bit(sys_rlreq) xor to_bit(sys_rlrdy))='0' then
				adjdqs_req <= to_stdulogic(to_bit(adjdqs_rdy));
				adjdqi_req <= to_stdulogic(to_bit(adjsto_rdy));
				adjsto_req <= to_stdulogic(to_bit(adjsto_rdy));
				state := sync_start;
			else
				case state is
				when sync_start =>
					if sys_sti(0)='1' then
						adjdqs_req <= not to_stdulogic(to_bit(adjdqs_rdy));
						state := sync_dqs;
					end if;
				when sync_dqs =>
					if (to_bit(adjdqs_req) xor to_bit(adjdqs_rdy))='0' then
						adjdqi_req <= not to_stdulogic(to_bit(adjsto_req));
						state := sync_dqi;
					end if;
				when sync_dqi =>
					if (adjsto_req xor adjdqi_req)='0' then
						adjsto_req <= not adjsto_rdy;
						state := sync_sto;
					end if;
				when sync_sto =>
					if (adjsto_req xor adjdqi_req)='0' then
						sys_rlrdy <= sys_rlreq;
						state := sync_start;
					end if;
				end case;

				aux := '1';
				for i in adjdqi_rdy'range loop
					aux := aux and (to_bit(adjdqi_rdy(i)) xor to_bit(adjdqi_req));
				end loop;
				adjsto_req <= to_stdulogic(aux) xor to_stdulogic(to_bit(adjdqi_req));
			end if;
		end if;
	end process;

	sys_rlcal <= to_stdulogic(to_bit(adjsto_req) xor to_bit(adjsto_rdy));

	dqsi_b : block
		signal step_rdy : std_logic;
		signal step_req : std_logic;
		signal delay    : std_logic_vector(0 to 5-1);
		signal dqsi     : std_logic;
		signal ddqsi    : std_logic;
		signal smp      : std_logic_vector(0 to DATA_GEAR-1);
		signal sto      : std_logic;
		signal imdr_rst : std_logic;
		signal imdr_clk : std_logic_vector(0 to 5-1);
	begin

		step_delay_e : entity hdl4fpga.align
		generic map (
			n => 1,
			d => (0 => 4))
		port map (
			clk => sys_clks(iodclk),
			di(0) => step_req,
			do(0) => step_rdy);

		adjdqs_e : entity hdl4fpga.adjpha
		generic map (
--			dtaps   => (taps+7)/8,
--			dtaps   => (taps+3)/4,
			taps    => taps)
		port map (
			edge     => std_logic'('1'),
			clk      => sys_clks(iodclk),
			req      => adjdqs_req,
			rdy      => adjdqs_rdy,
			step_req => step_req,
			step_rdy => step_rdy,
			smp      => smp,
			ph180    => dqs180,
			delay    => delay);

		ddqsi <= transport ddr_dqsi after dqs_linedelay;
		dqsidelay_i : idelaye2
		generic map (
			DELAY_SRC      => "IDATAIN",
			IDELAY_TYPE    => "VAR_LOAD",
			SIGNAL_PATTERN => "CLOCK")
		port map (
			regrst     => sys_rsts(rstiod),
			c          => sys_clks(iodclk),
			ld         => '1',
			cntvaluein => delay,
			idatain    => ddqsi,
			dataout    => dqsi_buf,
			cinvctrl   => '0',
			ce         => '0',
			inc        => '0',
			ldpipeen   => '0',
			datain     => '0');
			dqsi       <= dqsi_buf;

		imdr_clk <= (
			0 => sys_clks(clk0div),
			1 => sys_clks(clk0),
			2 => not sys_clks(clk90),
			3 => not sys_clks(clk0),
			4 => sys_clks(clk90));

		imdr_i : entity hdl4fpga.imdr
		generic map (
			SIZE => 1,
			GEAR => DATA_GEAR)
		port map (
			rst  => imdr_rst,
			clk  => imdr_clk,
			d(0) => dqsi,
			q    => smp);

		tp_dqsdly <= delay;
		process (sys_clks(clk0div))
		begin
			if rising_edge(sys_clks(clk0div)) then
				imdr_rst <= sys_rsts(rst0div);
			end if;
		end process;

		adjsto_e : entity hdl4fpga.adjsto
		generic map (
			GEAR => DATA_GEAR)
		port map (
			tp       => tp_dqssel,
			ddr_clk  => sys_clks(clk0div),
			edge     => '0',
			ddr_sti  => sys_sti(0),
			ddr_sto  => sto,
			dqs_smp  => smp,
			dqs_pre  => dqspre,
			sys_req  => adjsto_req,
			sys_rdy  => adjsto_rdy);

		process (sys_clks(clk90div))
			variable q : std_logic;
		begin
			if rising_edge(sys_clks(clk90div)) then
				if (not dqspre and dqs180)='1' then
					sys_sto <= (others => sto);
				elsif (not dqspre and not dqs180)='1' then
					sys_sto <= (others => sto);
				else
					sys_sto <= (others => q);
				end if;
				q := sto;
			end if;
		end process;

	end block;

	iod_rst <= not adjdqs_req;
	iddr_g : for i in ddr_dqi'range generate
		signal imdr_rst  : std_logic;
		signal imdr_clk  : std_logic_vector(0 to 5-1);
		signal adjdqi_st : std_logic;
	begin

		adjdqi_b : block
			signal delay    : std_logic_vector(0 to 5-1);
			signal step_req : std_logic;
			signal step_rdy : std_logic;
			signal dq_smp   : std_logic_vector(0 to DATA_GEAR-1);
			signal ddqi     : std_logic;
		begin

			step_delay_e : entity hdl4fpga.align
			generic map (
				n => 1,
				d => (0 => 4))
			port map (
				clk   => sys_clks(iodclk),
				di(0) => step_req,
				do(0) => step_rdy);

			dq_smp <= (dq(0*BYTE_SIZE+i), dq(1*BYTE_SIZE+i), dq(2*BYTE_SIZE+i), dq(3*BYTE_SIZE+i));
			adjdqi_e : entity hdl4fpga.adjpha
			generic map (
--				dtaps    => (taps+7)/8,
--				dtaps    => (taps+3)/4,
				taps     => taps)
			port map (
				edge     => std_logic'('0'),
				clk      => sys_clks(iodclk),
				req      => adjdqi_req,
				rdy      => adjdqi_rdy(i),
				step_req => step_req,
				step_rdy => step_rdy,
				smp      => dq_smp,
				delay    => delay);

			tp_g : if i=0 generate
				tp_dqidly <= delay;
			end generate;

			ddqi <= transport ddr_dqi(i) after dqi_linedelay;
			dqi_i : idelaye2
			generic map (
				DELAY_SRC    => "IDATAIN",
				IDELAY_TYPE  => "VAR_LOAD")
			port map (
				regrst      => iod_rst,
				c           => sys_clks(iodclk),
				ld          => '1',
				cntvaluein  => delay,
				idatain     => ddqi,
				dataout     => dqi(i),
				cinvctrl    => std_logic'('0'),
				ce          => std_logic'('0'),
				inc         => std_logic'('0'),
				ldpipeen    => std_logic'('0'),
				datain      => std_logic'('0'));

		end block;

		imdr_clk <= (
			0 => sys_clks(clk90div),
			1 => sys_clks(clk90),
			2 => sys_clks(clk90),
			3 => not sys_clks(clk90),
			4 => not sys_clks(clk90));

		process (sys_clks(clk90div))
			variable q : std_logic;
		begin
			if rising_edge(sys_clks(clk90div)) then
				imdr_rst <= q;
				q := sys_rsts(rst90div) or not adjdqs_req;
			end if;
		end process;

		imdr_i : entity hdl4fpga.imdr
		generic map (
			SIZE => 1,
			GEAR => DATA_GEAR)
		port map (
			rst  => imdr_rst,
			clk  => imdr_clk,
			d(0) => dqi(i),
			q(0) => dq(0*BYTE_SIZE+i),
			q(1) => dq(1*BYTE_SIZE+i),
			q(2) => dq(2*BYTE_SIZE+i),
			q(3) => dq(3*BYTE_SIZE+i));

		dly_b : block
		begin
			dly0_g : entity hdl4fpga.align
			generic map (
				n => 4,
				d => (0, 0, 1, 1))
			port map (
				clk => sys_clks(clk90div),
				di(0) => dq(0*BYTE_SIZE+i),
				di(1) => dq(1*BYTE_SIZE+i),
				di(2) => dq(2*BYTE_SIZE+i),
				di(3) => dq(3*BYTE_SIZE+i),
				do(0) => dqh(2*BYTE_SIZE+i),
				do(1) => dqh(3*BYTE_SIZE+i),
				do(2) => dqh(0*BYTE_SIZE+i),
				do(3) => dqh(1*BYTE_SIZE+i));

			dly1_g : entity hdl4fpga.align
			generic map (
				n => 4,
				d => (1, 1, 1, 1))
			port map (
				clk => sys_clks(clk90div),
				di(0) => dq(0*BYTE_SIZE+i),
				di(1) => dq(1*BYTE_SIZE+i),
				di(2) => dq(2*BYTE_SIZE+i),
				di(3) => dq(3*BYTE_SIZE+i),
				do(0) => dqf(0*BYTE_SIZE+i),
				do(1) => dqf(1*BYTE_SIZE+i),
				do(2) => dqf(2*BYTE_SIZE+i),
				do(3) => dqf(3*BYTE_SIZE+i));

		end block;

	end generate;
	sys_dqo <= dqh when (dqspre xor dqs180)='0' else dqf;

	oddr_g : for i in 0 to BYTE_SIZE-1 generate
		signal dqo   : std_logic_vector(0 to DATA_GEAR-1);
		signal clks  : std_logic_vector(0 to 2-1);
		signal dqt   : std_logic_vector(sys_dqt'range);
		signal dqclk : std_logic_vector(0 to 2-1);
		signal dq000 : std_logic_vector(0 to 2*DATA_GEAR-1);
		signal dq270 : std_logic_vector(0 to 2*DATA_GEAR-1);
		signal dq180 : std_logic_vector(0 to 2*DATA_GEAR-1);
		signal dq090 : std_logic_vector(0 to 2*DATA_GEAR-1);
	begin

		dqclk <= (0 => sys_clks(clk90div), 1 => sys_clks(clk90));

		clks <=
			(0 => sys_clks(clk90div), 1 => not sys_clks(clk90div)) when DATA_EDGE else
			(0 => sys_clks(clk90div), 1 => sys_clks(clk90div));

		registered_g : for j in clks'range generate
			gear_g : for l in 0 to DATA_GEAR/clks'length-1 generate
				process (sys_rlrdy, sys_rlreq, clks(j))
				begin
					if (to_bit(sys_rlrdy) xor to_bit(sys_rlreq))='1' then
						if j mod 2=1 then
							dqo(l*DATA_GEAR/clks'length+j) <= '1';
						else
							dqo(l*DATA_GEAR/clks'length+j) <= '0';
						end if;
					elsif rising_edge(clks(j)) then
						dqo(l*DATA_GEAR/clks'length+j) <= sys_dqi((l*DATA_GEAR/clks'length+j)*BYTE_SIZE+i);
					end if;
					if rising_edge(clks(j)) then
						dqt(l*DATA_GEAR/clks'length+j) <= reverse(sys_dqt)(l*DATA_GEAR/clks'length+j);
					end if;
				end process;
			end generate;
		end generate;

		omdr_i : entity hdl4fpga.omdr
		generic map (
			SIZE => 1,
			GEAR => DATA_GEAR)
		port map (
			rst   => sys_rsts(rst90div),
			clk   => dqclk,
			t     => dqt,
			tq(0) => ddr_dqt(i),
			d     => dqo,
			q(0)  => ddr_dqo(i));

	end generate;

	dmo_g : block
		signal dmt   : std_logic_vector(sys_dmt'range);
		signal dmi   : std_logic_vector(sys_dmi'range);
		signal clks  : std_logic_vector(0 to 2-1);
		signal dqclk : std_logic_vector(0 to 2-1);
		signal dq270 : std_logic_vector(0 to DATA_GEAR-1);
		signal dq180 : std_logic_vector(0 to DATA_GEAR-1);
		signal dq090 : std_logic_vector(0 to DATA_GEAR-1);
	begin

		dqclk <= (0 => sys_clks(clk90div), 1 => sys_clks(clk90));

		clks <=
			(0 => sys_clks(clk90div), 1 => not sys_clks(clk90div)) when DATA_EDGE else
			(0 => sys_clks(clk90div), 1 => sys_clks(clk90div));

		registered_g : for i in clks'range generate
			gear_g : for l in 0 to DATA_GEAR/clks'length-1 generate
				process (clks(i))
				begin
					if rising_edge(clks(i)) then
						dmi(l*DATA_GEAR/clks'length+i) <= sys_dmi(l*DATA_GEAR/clks'length+i);
					end if;
				end process;
			end generate;
		end generate;

		omdr_i : entity hdl4fpga.omdr
		generic map (
			SIZE => 1,
			GEAR => DATA_GEAR)
		port map (
			rst   => sys_rsts(rst90div),
			clk   => dqclk,
			t     => (others => '0'),
			tq(0) => ddr_dmt,
			d     => dmi,
			q(0)  => ddr_dmo);

	end block;

	dqso_b : block
		signal dqso      : std_logic_vector(sys_dqso'range);
		signal dqst      : std_logic_vector(sys_dqst'range);
		signal dqsclk    : std_logic_vector(0 to 2-1);
		signal adjdly    : std_logic_vector(0 to 5);
		signal adjdqs_st : std_logic;
	begin

		process (sys_dqso)
		begin
			dqso <= (others => '0');
			for i in dqso'range loop
				if i mod 2 = 1 then
					dqso(i) <= reverse(sys_dqso)(i);
				end if;
			end loop;
		end process;
		dqst <= reverse(sys_dqst);

		dqsclk <= (0 => sys_clks(clk0div), 1 => sys_clks(clk0));
		omdr_i : entity hdl4fpga.omdr
		generic map (
			SIZE => 1,
			GEAR => DATA_GEAR)
		port map (
			rst  => sys_rsts(rst0div),
			clk  => dqsclk,
			t    => dqst,
			tq(0)=> ddr_dqst,
			d    => dqso,
			q(0) => ddr_dqso);

	end block;
end;
