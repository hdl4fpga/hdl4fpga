library ieee;
use ieee.std_logic_1164.all;

package cgafonts6 is

	constant psf1digit8x8 : std_logic_vector(0 to 16*8*8-1) := (
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"00011000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"00000110" &
		B"01111100" &
		B"11000000" &
		B"11000000" &
		B"11111110" &
		B"00000000" &

		B"11111100" &
		B"00000110" &
		B"00000110" &
		B"00111100" &
		B"00000110" &
		B"00000110" &
		B"11111100" &
		B"00000000" &

		B"00001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11111110" &
		B"00001100" &
		B"00001100" &
		B"00000000" &

		B"11111110" &
		B"11000000" &
		B"11111100" &
		B"00000110" &
		B"00000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"01111100" &
		B"11000000" &
		B"11000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11111110" &
		B"00000110" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00110000" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"00000110" &
		B"01111100" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000"
		);

end;
