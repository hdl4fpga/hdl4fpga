-- (c) EMARD
-- License=BSD

library ieee;
use ieee.std_logic_1164.all;

package spi_display_init_pack is
  type T_spi_display_init_seq is array (natural range <>) of std_logic_vector(7 downto 0);
end;
