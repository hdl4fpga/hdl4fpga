--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library hdl4fpga;
use hdl4fpga.std.all;

entity sio_glue is
	port (
		sio_clk : in  std_logic;
		si_frm  : in  std_logic;
		si_irdy : in  std_logic;
		si_trdy : out std_logic;
		si_data : in  std_logic_vector;
		so_frm  : out std_logic;
		so_irdy : out std_logic;
		so_trdy : in  std_logic;
		so_data : out std_logic_vector);
end;

architecture def of sio_glue is
	signal des_data : std_logic_vector(0 to 8-1);
	signal ena : std_logic;
begin

	serdes_e : entity hdl4fpga.serdes
	port (
		serdes_clk => sio_clk
		serdes_frm => si_frm,
		ser_irdy   => si_irdy,
		ser_trdy   => open,
		ser_data   => si_data,

		des_frm    => des_frm,
		des_irdy   => des_irdy,
		des_data   => des_data);

	entity desser is
		port (
			desser_clk : in  std_logic;
	
			des_frm    : in  std_logic;
			des_irdy   : in  std_logic := '1';
			des_trdy   : out std_logic;
			des_data   : in  std_logic_vector;
	
			ser_irdy   : out std_logic;
			ser_trdy   : in  std_logic := '1';
			ser_data   : out std_logic_vector);
	end;

	process (sio_clk)
	begin
		if rising_edge(sio_clk) then
			if si_frm='0' then
				ena <= '0';
			elsif des_irdy='1' then
				ena <= '1';
			end if;
		end if;
	end process;

	tag_e : entity sio_tag is
	port map (
		sio_clk => sio_clk,
		sio_tag =>
		si_frm  => si_frm
		si_irdy : in  std_logic;
		si_trdy : out std_logic;
		si_data : in  std_logic_vector;
		so_frm  : out std_logic;
		so_irdy : out std_logic;
		so_trdy : in  std_logic;
		so_data : out std_logic_vector);

end;
