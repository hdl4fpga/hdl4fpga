package test is
	type std is ('0', '1');
end;

