library ieee;
use ieee.std_logic_1164.all;

package cgafonts1 is

	constant psf1bcd4x4 : std_logic_vector(0 to 16*4*4-1) := (
		B"1110" &
		B"1010" &
		B"1010" &
		B"1110" &

		B"0100" &
		B"1100" &
		B"0100" &
		B"1110" &

		B"1110" &
		B"0010" &
		B"1100" &
		B"1110" &
	
		B"1110" &
		B"0110" &
		B"0010" &
		B"1110" &
--	
		B"1010" &
		B"1110" &
		B"0010" &
		B"0010" &
	
		B"1100" &
		B"1110" &
		B"0010" &
		B"1110" &
	
		B"1000" &
		B"1110" &
		B"1010" &
		B"1110" &
	
		B"1110" &
		B"0010" &
		B"0100" &
		B"0100" &
--	
		B"1110" &
		B"1110" &
		B"1010" &
		B"1110" &
	
		B"1110" &
		B"1010" &
		B"1110" &
		B"0110" &
	
		B"0000" &
		B"0000" &
		B"0000" &
		B"0000" &

		B"0000" &
		B"0000" &
		B"0110" &
		B"0110" &
--		
		B"0100" &
		B"1110" &
		B"0100" &
		B"0000" &
	
		B"0000" &
		B"0110" &
		B"0000" &
		B"0000" &
	
		B"0000" &
		B"0000" &
		B"1111" &
		B"0000" &
	
		B"0000" &
		B"0000" &
		B"0000" &
		B"0000" );

end;