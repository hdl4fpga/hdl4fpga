library ieee;
use ieee.std_logic_1164.all
use ieee.numeric_std.all;

entity ecp3versa is
	port (
	);
end;

architecture scope of ecp3versa is
end;