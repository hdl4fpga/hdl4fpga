--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity imdr is
	generic (
		SIZE : natural;
		GEAR : natural);
	port (
		rst  : in  std_logic;
		clk  : in  std_logic_vector(0 to 5-1);
		ctrl : in  std_logic_vector(0 to 2-1) := (others => '0');
		d    : in  std_logic_vector(0 to SIZE-1);
		q    : out std_logic_vector(0 to SIZE*GEAR-1));
end;

library unisim;
use unisim.vcomponents.all;

architecture beh of imdr is
begin

	reg_g : for i in d'range generate
		signal po : std_logic_vector(0 to 4-1);
	begin

		iser_i : iserdese2
		generic map (
			INTERFACE_TYPE => "MEMORY",
			IOBDELAY => "BOTH",
			DYN_CLKDIV_INV_EN => "TRUE",
			DYN_CLK_INV_EN => "TRUE",
			NUM_CE => 1)
		port map (
			rst          => rst,
			dynclksel    => ctrl(1),
			clk          => clk(0),
			clkb         => clk(1),
			dynclkdivsel => ctrl(0),
			oclk         => clk(2),
			oclkb        => clk(3),
			clkdiv       => clk(4),
			ddly         => d(i),
			q1           => po(0),
			q2           => po(1),
			q3           => po(2),
			q4           => po(3),

			bitslip      => '0',
			ce1          => '1',
			ce2          => '1',
			clkdivp      => '0',
			d            => '0', --d(i),
			ofb          => '0',
			shiftin1     => '0',
			shiftin2     => '0');

		process (po)
		begin
			for j in 0 to GEAR-1 loop
				q(GEAR*i+j) <= po(j);
			end loop;
		end process;

	end generate;

end;
