library ieee;
use ieee.std_logic_1164.all;

package cgafonts5 is

	constant psf1cp850x8x8 : std_logic_vector(0 to 256*8*8-1) := (

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"01111110" &
		B"10000001" &
		B"10100101" &
		B"10000001" &
		B"10011101" &
		B"10111001" &
		B"10000001" &
		B"01111110" &

		B"01111110" &
		B"11111111" &
		B"11011011" &
		B"11111111" &
		B"11100011" &
		B"11000111" &
		B"11111111" &
		B"01111110" &

		B"01101100" &
		B"11111110" &
		B"11111110" &
		B"11111110" &
		B"01111100" &
		B"00111000" &
		B"00010000" &
		B"00000000" &

		B"00010000" &
		B"00111000" &
		B"01111100" &
		B"11111110" &
		B"01111100" &
		B"00111000" &
		B"00010000" &
		B"00000000" &

		B"00111000" &
		B"01111100" &
		B"00111000" &
		B"11111110" &
		B"11111110" &
		B"00010000" &
		B"00010000" &
		B"01111100" &

		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"11111111" &
		B"01111110" &
		B"00011000" &
		B"01111110" &

		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"00111100" &
		B"00011000" &
		B"00000000" &
		B"00000000" &

		B"11111111" &
		B"11111111" &
		B"11100111" &
		B"11000011" &
		B"11000011" &
		B"11100111" &
		B"11111111" &
		B"11111111" &

		B"00000000" &
		B"00111100" &
		B"01100110" &
		B"01000010" &
		B"01000010" &
		B"01100110" &
		B"00111100" &
		B"00000000" &

		B"11111111" &
		B"11000011" &
		B"10011001" &
		B"10111101" &
		B"10111101" &
		B"10011001" &
		B"11000011" &
		B"11111111" &

		B"00001111" &
		B"00000111" &
		B"00001111" &
		B"01111101" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"01111000" &

		B"00111100" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00011000" &
		B"01111110" &
		B"00011000" &

		B"00111111" &
		B"00110011" &
		B"00111111" &
		B"00110000" &
		B"00110000" &
		B"01110000" &
		B"11110000" &
		B"11100000" &

		B"01111111" &
		B"01100011" &
		B"01111111" &
		B"01100011" &
		B"01100011" &
		B"01100111" &
		B"11100110" &
		B"11000000" &

		B"10011001" &
		B"01011010" &
		B"00111100" &
		B"11100111" &
		B"11100111" &
		B"00111100" &
		B"01011010" &
		B"10011001" &

		B"10000000" &
		B"11100000" &
		B"11111000" &
		B"11111110" &
		B"11111000" &
		B"11100000" &
		B"10000000" &
		B"00000000" &

		B"00000010" &
		B"00001110" &
		B"00111110" &
		B"11111110" &
		B"00111110" &
		B"00001110" &
		B"00000010" &
		B"00000000" &

		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00111100" &
		B"00011000" &

		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00000000" &
		B"01100110" &
		B"00000000" &

		B"01111111" &
		B"11011011" &
		B"11011011" &
		B"01111011" &
		B"00011011" &
		B"00011011" &
		B"00011011" &
		B"00000000" &

		B"00111111" &
		B"01100000" &
		B"01111100" &
		B"01100110" &
		B"01100110" &
		B"00111110" &
		B"00000110" &
		B"11111100" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"01111110" &
		B"01111110" &
		B"00000000" &

		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"00011000" &
		B"01111110" &
		B"00111100" &
		B"00011000" &
		B"11111111" &

		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00111100" &
		B"00011000" &
		B"00000000" &

		B"00000000" &
		B"00011000" &
		B"00001100" &
		B"11111110" &
		B"00001100" &
		B"00011000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00110000" &
		B"01100000" &
		B"11111110" &
		B"01100000" &
		B"00110000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11111110" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00100100" &
		B"01100110" &
		B"11111111" &
		B"01100110" &
		B"00100100" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00011000" &
		B"00111100" &
		B"01111110" &
		B"11111111" &
		B"11111111" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"11111111" &
		B"11111111" &
		B"01111110" &
		B"00111100" &
		B"00011000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00011000" &
		B"00000000" &

		B"01101100" &
		B"01101100" &
		B"01101100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"01101100" &
		B"01101100" &
		B"11111110" &
		B"01101100" &
		B"11111110" &
		B"01101100" &
		B"01101100" &
		B"00000000" &

		B"00011000" &
		B"01111110" &
		B"11000000" &
		B"01111100" &
		B"00000110" &
		B"11111100" &
		B"00011000" &
		B"00000000" &

		B"00000000" &
		B"11000110" &
		B"11001100" &
		B"00011000" &
		B"00110000" &
		B"01100110" &
		B"11000110" &
		B"00000000" &

		B"00111000" &
		B"01101100" &
		B"00111000" &
		B"01110110" &
		B"11011100" &
		B"11001100" &
		B"01110110" &
		B"00000000" &

		B"00110000" &
		B"00110000" &
		B"01100000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00000000" &

		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00000000" &

		B"00000000" &
		B"01100110" &
		B"00111100" &
		B"11111111" &
		B"00111100" &
		B"01100110" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00110000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11000000" &
		B"10000000" &
		B"00000000" &

		B"01111100" &
		B"11001110" &
		B"11011110" &
		B"11110110" &
		B"11100110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"00011000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"00000110" &
		B"01111100" &
		B"11000000" &
		B"11000000" &
		B"11111110" &
		B"00000000" &

		B"11111100" &
		B"00000110" &
		B"00000110" &
		B"00111100" &
		B"00000110" &
		B"00000110" &
		B"11111100" &
		B"00000000" &

		B"00001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11111110" &
		B"00001100" &
		B"00001100" &
		B"00000000" &

		B"11111110" &
		B"11000000" &
		B"11111100" &
		B"00000110" &
		B"00000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"01111100" &
		B"11000000" &
		B"11000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11111110" &
		B"00000110" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00110000" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"00000110" &
		B"01111100" &
		B"00000000" &

		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00110000" &

		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"00000000" &

		B"00111100" &
		B"01100110" &
		B"00001100" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00011000" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11011110" &
		B"11011110" &
		B"11011110" &
		B"11000000" &
		B"01111110" &
		B"00000000" &

		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11111100" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11111000" &
		B"11001100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11001100" &
		B"11111000" &
		B"00000000" &

		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11111000" &
		B"11000000" &
		B"11000000" &
		B"11111110" &
		B"00000000" &

		B"11111110" &
		B"11000000" &
		B"11000000" &
		B"11111000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"11000000" &
		B"11001110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00000000" &

		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11000110" &
		B"11001100" &
		B"11011000" &
		B"11110000" &
		B"11011000" &
		B"11001100" &
		B"11000110" &
		B"00000000" &

		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11111110" &
		B"00000000" &

		B"11000110" &
		B"11101110" &
		B"11111110" &
		B"11111110" &
		B"11010110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"11000110" &
		B"11100110" &
		B"11110110" &
		B"11011110" &
		B"11001110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11111100" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11010110" &
		B"11011110" &
		B"01111100" &
		B"00000110" &

		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11111100" &
		B"11011000" &
		B"11001100" &
		B"11000110" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"01111100" &
		B"00000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11111111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"00000000" &

		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00111000" &
		B"00000000" &

		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11010110" &
		B"11111110" &
		B"01101100" &
		B"00000000" &

		B"11000110" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00011000" &
		B"00110000" &
		B"11100000" &
		B"00000000" &

		B"11111110" &
		B"00000110" &
		B"00001100" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11111110" &
		B"00000000" &

		B"00111100" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00110000" &
		B"00111100" &
		B"00000000" &

		B"11000000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00001100" &
		B"00000110" &
		B"00000010" &
		B"00000000" &

		B"00111100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"00111100" &
		B"00000000" &

		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &

		B"00011000" &
		B"00011000" &
		B"00001100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"00000110" &
		B"01111110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11111100" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"01111110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"01111100" &
		B"00000000" &

		B"00011100" &
		B"00110110" &
		B"00110000" &
		B"01111000" &
		B"00110000" &
		B"00110000" &
		B"01111000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"11111100" &

		B"11000000" &
		B"11000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"00011000" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &

		B"00000110" &
		B"00000000" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"00000110" &
		B"11000110" &
		B"01111100" &

		B"11000000" &
		B"11000000" &
		B"11001100" &
		B"11011000" &
		B"11111000" &
		B"11001100" &
		B"11000110" &
		B"00000000" &

		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11001100" &
		B"11111110" &
		B"11111110" &
		B"11010110" &
		B"11010110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11111100" &
		B"11000000" &
		B"11000000" &

		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"00000110" &

		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"11000110" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"11000000" &
		B"01111100" &
		B"00000110" &
		B"11111100" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00001110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00111000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11010110" &
		B"11111110" &
		B"01101100" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"01101100" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000110" &
		B"11111100" &

		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"00001100" &
		B"00111000" &
		B"01100000" &
		B"11111110" &
		B"00000000" &

		B"00001110" &
		B"00011000" &
		B"00011000" &
		B"01110000" &
		B"00011000" &
		B"00011000" &
		B"00001110" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"01110000" &
		B"00011000" &
		B"00011000" &
		B"00001110" &
		B"00011000" &
		B"00011000" &
		B"01110000" &
		B"00000000" &

		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00010000" &
		B"00111000" &
		B"01101100" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"00000000" &

		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11010110" &
		B"01111100" &
		B"00110000" &

		B"11000110" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"00001110" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"01111100" &
		B"00000000" &

		B"01111110" &
		B"10000001" &
		B"00111100" &
		B"00000110" &
		B"01111110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"01100110" &
		B"00000000" &
		B"01111100" &
		B"00000110" &
		B"01111110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"11100000" &
		B"00000000" &
		B"01111100" &
		B"00000110" &
		B"01111110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"01111100" &
		B"00000110" &
		B"01111110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000000" &
		B"11010110" &
		B"01111100" &
		B"00110000" &

		B"01111110" &
		B"10000001" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"01111100" &
		B"00000000" &

		B"01100110" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"01111100" &
		B"00000000" &

		B"11100000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000000" &
		B"01111100" &
		B"00000000" &

		B"01100110" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &

		B"01111100" &
		B"10000010" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &

		B"01110000" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &

		B"11000110" &
		B"00010000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"00111000" &
		B"00111000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11111110" &
		B"11000110" &
		B"00000000" &

		B"00001110" &
		B"00000000" &
		B"11111110" &
		B"11000000" &
		B"11111000" &
		B"11000000" &
		B"11111110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111111" &
		B"00001100" &
		B"01111111" &
		B"11001100" &
		B"01111111" &
		B"00000000" &

		B"00111111" &
		B"01101100" &
		B"11001100" &
		B"11111111" &
		B"11001100" &
		B"11001100" &
		B"11001111" &
		B"00000000" &

		B"01111100" &
		B"10000010" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"01100110" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11100000" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"01111100" &
		B"10000010" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"11100000" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"01100110" &
		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"00111110" &
		B"00000110" &
		B"01111100" &

		B"11000110" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"11000110" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11111110" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"11011000" &
		B"11011000" &
		B"11011000" &
		B"01111110" &
		B"00011000" &

		B"00111000" &
		B"01101100" &
		B"01100000" &
		B"11110000" &
		B"01100000" &
		B"01100110" &
		B"11111100" &
		B"00000000" &

		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"01111110" &
		B"00011000" &

		B"11111000" &
		B"11001100" &
		B"11001100" &
		B"11111010" &
		B"11000110" &
		B"11001111" &
		B"11000110" &
		B"11000011" &

		B"00001110" &
		B"00011011" &
		B"00011000" &
		B"00111100" &
		B"00011000" &
		B"00011000" &
		B"11011000" &
		B"01110000" &

		B"00001110" &
		B"00000000" &
		B"01111100" &
		B"00000110" &
		B"01111110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"00011100" &
		B"00000000" &
		B"00111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00111100" &
		B"00000000" &

		B"00001110" &
		B"00000000" &
		B"01111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"00001110" &
		B"00000000" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"01111110" &
		B"00000000" &

		B"00000000" &
		B"11111110" &
		B"00000000" &
		B"11111100" &
		B"11000110" &
		B"11000110" &
		B"11000110" &
		B"00000000" &

		B"11111110" &
		B"00000000" &
		B"11000110" &
		B"11100110" &
		B"11110110" &
		B"11011110" &
		B"11001110" &
		B"00000000" &

		B"00111100" &
		B"01101100" &
		B"01101100" &
		B"00111110" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &

		B"00111100" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &

		B"00011000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00110000" &
		B"01100110" &
		B"00111100" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"11000000" &
		B"11000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111100" &
		B"00001100" &
		B"00001100" &
		B"00000000" &
		B"00000000" &

		B"11000110" &
		B"11001100" &
		B"11011000" &
		B"00111111" &
		B"01100011" &
		B"11001111" &
		B"10001100" &
		B"00001111" &

		B"11000011" &
		B"11000110" &
		B"11001100" &
		B"11011011" &
		B"00110111" &
		B"01101101" &
		B"11001111" &
		B"00000011" &

		B"00011000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"00000000" &
		B"00110011" &
		B"01100110" &
		B"11001100" &
		B"01100110" &
		B"00110011" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"11001100" &
		B"01100110" &
		B"00110011" &
		B"01100110" &
		B"11001100" &
		B"00000000" &
		B"00000000" &

		B"00100010" &
		B"10001000" &
		B"00100010" &
		B"10001000" &
		B"00100010" &
		B"10001000" &
		B"00100010" &
		B"10001000" &

		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &
		B"01010101" &
		B"10101010" &

		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &
		B"11011101" &
		B"01110111" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00011000" &
		B"00011000" &
		B"11111000" &
		B"00011000" &
		B"11111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"11110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00000000" &
		B"00000000" &
		B"11111000" &
		B"00011000" &
		B"11111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00110110" &
		B"00110110" &
		B"11110110" &
		B"00000110" &
		B"11110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"00000110" &
		B"11110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00110110" &
		B"00110110" &
		B"11110110" &
		B"00000110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"11111110" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"11111000" &
		B"00011000" &
		B"11111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11111111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00011000" &
		B"00011000" &
		B"00011111" &
		B"00011000" &
		B"00011111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00110110" &
		B"00110110" &
		B"00110111" &
		B"00110000" &
		B"00111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00111111" &
		B"00110000" &
		B"00110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00110110" &
		B"00110110" &
		B"11110111" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"11110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00110110" &
		B"00110110" &
		B"00110111" &
		B"00110000" &
		B"00110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00110110" &
		B"00110110" &
		B"11110111" &
		B"00000000" &
		B"11110111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00011000" &
		B"00011000" &
		B"11111111" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00000000" &
		B"11111111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"00011111" &
		B"00011000" &
		B"00011111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00011111" &
		B"00011000" &
		B"00011111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00111111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"00110110" &
		B"11111111" &
		B"00110110" &
		B"00110110" &
		B"00110110" &

		B"00011000" &
		B"00011000" &
		B"11111111" &
		B"00011000" &
		B"11111111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011111" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &

		B"11110000" &
		B"11110000" &
		B"11110000" &
		B"11110000" &
		B"11110000" &
		B"11110000" &
		B"11110000" &
		B"11110000" &

		B"00001111" &
		B"00001111" &
		B"00001111" &
		B"00001111" &
		B"00001111" &
		B"00001111" &
		B"00001111" &
		B"00001111" &

		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"11111111" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01110110" &
		B"11011100" &
		B"11001000" &
		B"11011100" &
		B"01110110" &
		B"00000000" &

		B"00111000" &
		B"01101100" &
		B"01101100" &
		B"01111000" &
		B"01101100" &
		B"01100110" &
		B"01101100" &
		B"01100000" &

		B"00000000" &
		B"11111110" &
		B"11000110" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"11000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"11111110" &
		B"01101100" &
		B"01101100" &
		B"01101100" &
		B"01101100" &
		B"00000000" &

		B"11111110" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"11111110" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"11011000" &
		B"11011000" &
		B"11011000" &
		B"01110000" &
		B"00000000" &

		B"00000000" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01100110" &
		B"01111100" &
		B"01100000" &
		B"11000000" &

		B"00000000" &
		B"01110110" &
		B"11011100" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"01111110" &
		B"00011000" &
		B"00111100" &
		B"01100110" &
		B"01100110" &
		B"00111100" &
		B"00011000" &
		B"01111110" &

		B"00111100" &
		B"01100110" &
		B"11000011" &
		B"11111111" &
		B"11000011" &
		B"01100110" &
		B"00111100" &
		B"00000000" &

		B"00111100" &
		B"01100110" &
		B"11000011" &
		B"11000011" &
		B"01100110" &
		B"01100110" &
		B"11100111" &
		B"00000000" &

		B"00001110" &
		B"00011000" &
		B"00001100" &
		B"01111110" &
		B"11000110" &
		B"11000110" &
		B"01111100" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"01111110" &
		B"11011011" &
		B"11011011" &
		B"01111110" &
		B"00000000" &
		B"00000000" &

		B"00000110" &
		B"00001100" &
		B"01111110" &
		B"11011011" &
		B"11011011" &
		B"01111110" &
		B"01100000" &
		B"11000000" &

		B"00111000" &
		B"01100000" &
		B"11000000" &
		B"11111000" &
		B"11000000" &
		B"01100000" &
		B"00111000" &
		B"00000000" &

		B"01111000" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"11001100" &
		B"00000000" &

		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00000000" &

		B"00011000" &
		B"00011000" &
		B"01111110" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"01111110" &
		B"00000000" &

		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"00000000" &
		B"11111100" &
		B"00000000" &

		B"00011000" &
		B"00110000" &
		B"01100000" &
		B"00110000" &
		B"00011000" &
		B"00000000" &
		B"11111100" &
		B"00000000" &

		B"00001110" &
		B"00011011" &
		B"00011011" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &

		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"00011000" &
		B"11011000" &
		B"11011000" &
		B"01110000" &

		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"01111110" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &

		B"00000000" &
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"01110110" &
		B"11011100" &
		B"00000000" &
		B"00000000" &

		B"00111000" &
		B"01101100" &
		B"01101100" &
		B"00111000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00011000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00001111" &
		B"00001100" &
		B"00001100" &
		B"00001100" &
		B"11101100" &
		B"01101100" &
		B"00111100" &
		B"00011100" &

		B"01111000" &
		B"01101100" &
		B"01101100" &
		B"01101100" &
		B"01101100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"01111100" &
		B"00001100" &
		B"01111100" &
		B"01100000" &
		B"01111100" &
		B"00000000" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00000000" &
		B"00111100" &
		B"00111100" &
		B"00111100" &
		B"00111100" &
		B"00000000" &
		B"00000000" &

		B"00000000" &
		B"00010000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000" &
		B"00000000"
		);

end;