--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

library ieee;
use ieee.std_logic_1164.all;

package cp850x8x8x0to127 is

	constant psf1cp850x8x8x0to127 : std_logic_vector(0*8*8 to 128*8*8-1) := (

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"01111110" &
		"10000001" &
		"10100101" &
		"10000001" &
		"10011101" &
		"10111001" &
		"10000001" &
		"01111110" &

		"01111110" &
		"11111111" &
		"11011011" &
		"11111111" &
		"11100011" &
		"11000111" &
		"11111111" &
		"01111110" &

		"01101100" &
		"11111110" &
		"11111110" &
		"11111110" &
		"01111100" &
		"00111000" &
		"00010000" &
		"00000000" &

		"00010000" &
		"00111000" &
		"01111100" &
		"11111110" &
		"01111100" &
		"00111000" &
		"00010000" &
		"00000000" &

		"00111000" &
		"01111100" &
		"00111000" &
		"11111110" &
		"11111110" &
		"00010000" &
		"00010000" &
		"01111100" &

		"00000000" &
		"00011000" &
		"00111100" &
		"01111110" &
		"11111111" &
		"01111110" &
		"00011000" &
		"01111110" &

		"00000000" &
		"00000000" &
		"00011000" &
		"00111100" &
		"00111100" &
		"00011000" &
		"00000000" &
		"00000000" &

		"11111111" &
		"11111111" &
		"11100111" &
		"11000011" &
		"11000011" &
		"11100111" &
		"11111111" &
		"11111111" &

		"00000000" &
		"00111100" &
		"01100110" &
		"01000010" &
		"01000010" &
		"01100110" &
		"00111100" &
		"00000000" &

		"11111111" &
		"11000011" &
		"10011001" &
		"10111101" &
		"10111101" &
		"10011001" &
		"11000011" &
		"11111111" &

		"00001111" &
		"00000111" &
		"00001111" &
		"01111101" &
		"11001100" &
		"11001100" &
		"11001100" &
		"01111000" &

		"00111100" &
		"01100110" &
		"01100110" &
		"01100110" &
		"00111100" &
		"00011000" &
		"01111110" &
		"00011000" &

		"00111111" &
		"00110011" &
		"00111111" &
		"00110000" &
		"00110000" &
		"01110000" &
		"11110000" &
		"11100000" &

		"01111111" &
		"01100011" &
		"01111111" &
		"01100011" &
		"01100011" &
		"01100111" &
		"11100110" &
		"11000000" &

		"10011001" &
		"01011010" &
		"00111100" &
		"11100111" &
		"11100111" &
		"00111100" &
		"01011010" &
		"10011001" &

		"10000000" &
		"11100000" &
		"11111000" &
		"11111110" &
		"11111000" &
		"11100000" &
		"10000000" &
		"00000000" &

		"00000010" &
		"00001110" &
		"00111110" &
		"11111110" &
		"00111110" &
		"00001110" &
		"00000010" &
		"00000000" &

		"00011000" &
		"00111100" &
		"01111110" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00111100" &
		"00011000" &

		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"01100110" &
		"00000000" &
		"01100110" &
		"00000000" &

		"01111111" &
		"11011011" &
		"11011011" &
		"01111011" &
		"00011011" &
		"00011011" &
		"00011011" &
		"00000000" &

		"00111111" &
		"01100000" &
		"01111100" &
		"01100110" &
		"01100110" &
		"00111110" &
		"00000110" &
		"11111100" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"01111110" &
		"01111110" &
		"01111110" &
		"00000000" &

		"00011000" &
		"00111100" &
		"01111110" &
		"00011000" &
		"01111110" &
		"00111100" &
		"00011000" &
		"11111111" &

		"00011000" &
		"00111100" &
		"01111110" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00111100" &
		"00011000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00001100" &
		"11111110" &
		"00001100" &
		"00011000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00110000" &
		"01100000" &
		"11111110" &
		"01100000" &
		"00110000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00100100" &
		"01100110" &
		"11111111" &
		"01100110" &
		"00100100" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00111100" &
		"01111110" &
		"11111111" &
		"11111111" &
		"00000000" &
		"00000000" &

		"00000000" &
		"11111111" &
		"11111111" &
		"01111110" &
		"00111100" &
		"00011000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00011000" &
		"00000000" &

		"01101100" &
		"01101100" &
		"01101100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"01101100" &
		"01101100" &
		"11111110" &
		"01101100" &
		"11111110" &
		"01101100" &
		"01101100" &
		"00000000" &

		"00011000" &
		"01111110" &
		"11000000" &
		"01111100" &
		"00000110" &
		"11111100" &
		"00011000" &
		"00000000" &

		"00000000" &
		"11000110" &
		"11001100" &
		"00011000" &
		"00110000" &
		"01100110" &
		"11000110" &
		"00000000" &

		"00111000" &
		"01101100" &
		"00111000" &
		"01110110" &
		"11011100" &
		"11001100" &
		"01110110" &
		"00000000" &

		"00110000" &
		"00110000" &
		"01100000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00001100" &
		"00011000" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00011000" &
		"00001100" &
		"00000000" &

		"00110000" &
		"00011000" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00011000" &
		"00110000" &
		"00000000" &

		"00000000" &
		"01100110" &
		"00111100" &
		"11111111" &
		"00111100" &
		"01100110" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00110000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"01111110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"01100000" &
		"11000000" &
		"10000000" &
		"00000000" &

		"01111100" &
		"11001110" &
		"11011110" &
		"11110110" &
		"11100110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00011000" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00000000" &

		"01111100" &
		"11000110" &
		"00000110" &
		"01111100" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &

		"11111100" &
		"00000110" &
		"00000110" &
		"00111100" &
		"00000110" &
		"00000110" &
		"11111100" &
		"00000000" &

		"00001100" &
		"11001100" &
		"11001100" &
		"11001100" &
		"11111110" &
		"00001100" &
		"00001100" &
		"00000000" &

		"11111110" &
		"11000000" &
		"11111100" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"01111100" &
		"11000000" &
		"11000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111110" &
		"00000110" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"00110000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"00000110" &
		"01111100" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"00000000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00110000" &

		"00001100" &
		"00011000" &
		"00110000" &
		"01100000" &
		"00110000" &
		"00011000" &
		"00001100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"00000000" &
		"01111110" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00110000" &
		"00011000" &
		"00001100" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"00000000" &

		"00111100" &
		"01100110" &
		"00001100" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00011000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11011110" &
		"11011110" &
		"11011110" &
		"11000000" &
		"01111110" &
		"00000000" &

		"00111000" &
		"01101100" &
		"11000110" &
		"11000110" &
		"11111110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111000" &
		"11001100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11001100" &
		"11111000" &
		"00000000" &

		"11111110" &
		"11000000" &
		"11000000" &
		"11111000" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &

		"11111110" &
		"11000000" &
		"11000000" &
		"11111000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000000" &
		"11000000" &
		"11001110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"11111110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"01111110" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"01111110" &
		"00000000" &

		"00000110" &
		"00000110" &
		"00000110" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11000110" &
		"11001100" &
		"11011000" &
		"11110000" &
		"11011000" &
		"11001100" &
		"11000110" &
		"00000000" &

		"11000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11000000" &
		"11111110" &
		"00000000" &

		"11000110" &
		"11101110" &
		"11111110" &
		"11111110" &
		"11010110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"11000110" &
		"11100110" &
		"11110110" &
		"11011110" &
		"11001110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"11000000" &
		"11000000" &
		"11000000" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11010110" &
		"11011110" &
		"01111100" &
		"00000110" &

		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"11011000" &
		"11001100" &
		"11000110" &
		"00000000" &

		"01111100" &
		"11000110" &
		"11000000" &
		"01111100" &
		"00000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"11111111" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11111110" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00111000" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11010110" &
		"11111110" &
		"01101100" &
		"00000000" &

		"11000110" &
		"11000110" &
		"01101100" &
		"00111000" &
		"01101100" &
		"11000110" &
		"11000110" &
		"00000000" &

		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00011000" &
		"00110000" &
		"11100000" &
		"00000000" &

		"11111110" &
		"00000110" &
		"00001100" &
		"00011000" &
		"00110000" &
		"01100000" &
		"11111110" &
		"00000000" &

		"00111100" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00110000" &
		"00111100" &
		"00000000" &

		"11000000" &
		"01100000" &
		"00110000" &
		"00011000" &
		"00001100" &
		"00000110" &
		"00000010" &
		"00000000" &

		"00111100" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00001100" &
		"00111100" &
		"00000000" &

		"00010000" &
		"00111000" &
		"01101100" &
		"11000110" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"11111111" &

		"00011000" &
		"00011000" &
		"00001100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"00000110" &
		"01111110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"11000000" &
		"11000000" &
		"11000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000000" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00000110" &
		"00000110" &
		"00000110" &
		"01111110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11111110" &
		"11000000" &
		"01111100" &
		"00000000" &

		"00011100" &
		"00110110" &
		"00110000" &
		"01111000" &
		"00110000" &
		"00110000" &
		"01111000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"11111100" &

		"11000000" &
		"11000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"00011000" &
		"00000000" &
		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00111100" &
		"00000000" &

		"00000110" &
		"00000000" &
		"00000110" &
		"00000110" &
		"00000110" &
		"00000110" &
		"11000110" &
		"01111100" &

		"11000000" &
		"11000000" &
		"11001100" &
		"11011000" &
		"11111000" &
		"11001100" &
		"11000110" &
		"00000000" &

		"00111000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11001100" &
		"11111110" &
		"11111110" &
		"11010110" &
		"11010110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111100" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11111100" &
		"11000110" &
		"11000110" &
		"11111100" &
		"11000000" &
		"11000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"00000110" &

		"00000000" &
		"00000000" &
		"11111100" &
		"11000110" &
		"11000000" &
		"11000000" &
		"11000000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"01111110" &
		"11000000" &
		"01111100" &
		"00000110" &
		"11111100" &
		"00000000" &

		"00011000" &
		"00011000" &
		"01111110" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00001110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111100" &
		"00111000" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11010110" &
		"11111110" &
		"01101100" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"01101100" &
		"00111000" &
		"01101100" &
		"11000110" &
		"00000000" &

		"00000000" &
		"00000000" &
		"11000110" &
		"11000110" &
		"11000110" &
		"01111110" &
		"00000110" &
		"11111100" &

		"00000000" &
		"00000000" &
		"11111110" &
		"00001100" &
		"00111000" &
		"01100000" &
		"11111110" &
		"00000000" &

		"00001110" &
		"00011000" &
		"00011000" &
		"01110000" &
		"00011000" &
		"00011000" &
		"00001110" &
		"00000000" &

		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &
		"00011000" &
		"00011000" &
		"00011000" &
		"00000000" &

		"01110000" &
		"00011000" &
		"00011000" &
		"00001110" &
		"00011000" &
		"00011000" &
		"01110000" &
		"00000000" &

		"01110110" &
		"11011100" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &
		"00000000" &

		"00000000" &
		"00010000" &
		"00111000" &
		"01101100" &
		"11000110" &
		"11000110" &
		"11111110" &
		"00000000");

end;

