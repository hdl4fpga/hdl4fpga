--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library hdl4fpga;
use hdl4fpga.std.all;

entity sio_hdlc is
	generic (
		mem_size  : natural := 4*(2048*8));
	port (
		uart_clk    : in  std_logic;

		uartrx_irdy : in  std_logic;
		uartrx_data : in  std_logic_vector;

		uarttx_irdy : out std_logic;
		uarttx_trdy : in  std_logic;
		uarttx_data : out std_logic_vector;

		sio_clk   : in  std_logic;
		si_frm    : in  std_logic;
		si_irdy   : in  std_logic;
		si_trdy   : buffer std_logic;
		si_end    : in  std_logic;
		si_data   : in  std_logic_vector;

		so_frm    : buffer std_logic;
		so_irdy   : out std_logic;
		so_trdy   : in  std_logic;
		so_data   : out std_logic_vector;
		tp : out std_logic_vector(1 to 32));
end;

architecture def of sio_hdlc is

	signal rx_frm  : std_logic;
	signal rx_irdy : std_logic;
	signal rx_trdy : std_logic;
	signal rx_end  : std_logic;
	signal rx_data : std_logic_vector(si_data'range);

	signal tx_frm  : std_logic;
	signal tx_irdy : std_logic;
	signal tx_trdy : std_logic;
	signal tx_data : std_logic_vector(si_data'range);

begin

	hdlc_b : block

		signal hdlcrx_frm    : std_logic;
		signal hdlcrx_irdy   : std_logic;
		signal hdlcrx_data   : std_logic_vector(so_data'range);

		signal hdlcfcsrx_sb  : std_logic;
		signal hdlcfcsrx_vld : std_logic;

		signal fifo_cmmt     : std_logic;
		signal fifo_avail    : std_logic;
		signal fifo_rllbk    : std_logic;

	begin

		hdlcdll_rx_e : entity hdl4fpga.hdlcdll_rx
		port map (
			uart_clk    => uart_clk,
			uartrx_irdy => uartrx_irdy,
			uartrx_data => uartrx_data,

			hdlcrx_frm  => hdlcrx_frm,
			hdlcrx_irdy => hdlcrx_irdy,
			hdlcrx_data => hdlcrx_data,
			fcs_sb      => hdlcfcsrx_sb,
			fcs_vld     => hdlcfcsrx_vld);

		fifo_cmmt  <= hdlcfcsrx_sb and     hdlcfcsrx_vld;
		fifo_rllbk <= hdlcfcsrx_sb and not hdlcfcsrx_vld;

		fifo_e : entity hdl4fpga.txn_buffer
		generic map (
			m => 11)
		port map (
			src_clk  => uart_clk,
			src_frm  => hdlcrx_frm,
			src_irdy => hdlcrx_irdy,
			src_trdy => open,
			src_data => hdlcrx_data,

			rollback => fifo_rllbk,
			commit   => fifo_cmmt,
			avail    => fifo_avail,

			dst_frm  => rx_frm,
			dst_irdy => rx_irdy,
			dst_trdy => rx_trdy,
			dst_end  => rx_end,
			dst_data => rx_data);

		rx_frm_p : process (sio_clk)
		begin
			if rising_edge(sio_clk) then
				if rx_frm='0' then
					if fifo_avail='1' then
						rx_frm <= '1';
					end if;
				elsif rx_end='1' and rx_trdy='1' then
					rx_frm <= '0';
				end if;
			end if;
		end process;

		rx_irdy <=
			'0'     when rx_frm='0' else
			rx_trdy when rx_end='0' else
			'0';

		hdlcdll_tx_e : entity hdl4fpga.hdlcdll_tx
		port map (
			uart_clk    => uart_clk,
			uart_irdy   => uarttx_irdy,
			uart_trdy   => uarttx_trdy,
			uart_data   => uarttx_data,

			hdlctx_frm  => si_frm,
			hdlctx_irdy => si_irdy,
			hdlctx_trdy => si_trdy,
			hdlctx_end  => si_end,
			hdlctx_data => si_data);

	end block;

	flow_e : entity hdl4fpga.sio_flow
	port map (
		tp      => tp,
		sio_clk => uart_clk,

		rx_frm  => rx_frm,
		rx_irdy => rx_irdy,
		rx_trdy => rx_trdy,
		rx_data => rx_data,

		so_frm  => so_frm,
		so_irdy => so_irdy,
		so_trdy => so_trdy,
		so_data => so_data,

		si_frm  => si_frm,
		si_irdy => si_irdy,
		si_trdy => si_trdy,
		si_data => si_data,

		tx_frm  => tx_frm,
		tx_irdy => tx_irdy,
		tx_trdy => tx_trdy,
		tx_data => tx_data);

end;
