--                                                                            --
-- Author(s):                                                                 --
--   Miguel Angel Sagreras                                                    --
--                                                                            --
-- Copyright (C) 2015                                                         --
--    Miguel Angel Sagreras                                                   --
--                                                                            --
-- This source file may be used and distributed without restriction provided  --
-- that this copyright statement is not removed from the file and that any    --
-- derivative work contains  the original copyright notice and the associated --
-- disclaimer.                                                                --
--                                                                            --
-- This source file is free software; you can redistribute it and/or modify   --
-- it under the terms of the GNU General Public License as published by the   --
-- Free Software Foundation, either version 3 of the License, or (at your     --
-- option) any later version.                                                 --
--                                                                            --
-- This source is distributed in the hope that it will be useful, but WITHOUT --
-- ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or      --
-- FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License for   --
-- more details at http://www.gnu.org/licenses/.                              --
--                                                                            --

library hdl4fpga;
use hdl4fpga.std.all;

architecture ulx3s_graphics of testbench is

	constant bank_bits  : natural := 2;
	constant addr_bits  : natural := 13;
	constant cols_bits  : natural := 9;
	constant data_bytes : natural := 2;
	constant byte_bits  : natural := 8;
	constant data_bits  : natural := byte_bits*data_bytes;

	signal rst   : std_logic;
	signal xtal  : std_logic := '0';

	signal sdram_dq    : std_logic_vector (data_bits - 1 downto 0) := (others => 'Z');
	signal sdram_addr  : std_logic_vector (addr_bits - 1 downto 0);
	signal sdram_ba    : std_logic_vector (1 downto 0);
	signal sdram_clk   : std_logic := '0';
	signal sdram_cke   : std_logic := '1';
	signal sdram_cs_n  : std_logic := '1';
	signal sdram_ras_n : std_logic;
	signal sdram_cas_n : std_logic;
	signal sdram_we_n  : std_logic;
	signal sdram_dqm   : std_logic_vector(1 downto 0);

	component ulx3s is
		port (
			clk_25mhz      : in    std_logic;

			ftdi_rxd       : out   std_logic;
			ftdi_txd       : in    std_logic := '-';
			ftdi_nrts      : inout std_logic := '-';
			ftdi_ndtr      : inout std_logic := '-';
			ftdi_txden     : inout std_logic := '-';

			led            : out   std_logic_vector(8-1 downto 0);
			btn            : in    std_logic_vector(7-1 downto 0) := (others => '-');
			sw             : in    std_logic_vector(4-1 downto 0) := (others => '-');


			oled_clk       : out   std_logic;
			oled_mosi      : out   std_logic;
			oled_dc        : out   std_logic;
			oled_resn      : out   std_logic;
			oled_csn       : out   std_logic;

			--flash_csn      : out   std_logic;
			--flash_clk      : out   std_logic;
			--flash_mosi     : out   std_logic;
			--flash_miso     : in    std_logic;
			--flash_holdn    : out   std_logic;
			--flash_wpn      : out   std_logic;

			sd_clk         : in    std_logic := '-';
			sd_cmd         : out   std_logic; -- sd_cmd=MOSI (out)
			sd_d           : inout std_logic_vector(4-1 downto 0) := (others => '-'); -- sd_d(0)=MISO (in), sd_d(3)=CSn (out)
			sd_wp          : in    std_logic := '-';
			sd_cdn         : in    std_logic := '-'; -- card detect not connected

			adc_csn        : out   std_logic;
			adc_mosi       : out   std_logic;
			adc_miso       : in    std_logic := '-';
			adc_sclk       : out   std_logic;

			audio_l        : out   std_logic_vector(4-1 downto 0);
			audio_r        : out   std_logic_vector(4-1 downto 0);
			audio_v        : out   std_logic_vector(4-1 downto 0);

			wifi_en        : out   std_logic := '1'; -- '0' disables ESP32
			wifi_rxd       : out   std_logic;
			wifi_txd       : in    std_logic := '-';
			wifi_gpio0     : out   std_logic := '1'; -- '0' requests ESP32 to upload "passthru" bitstream
			wifi_gpio5     : inout std_logic := '-';
			wifi_gpio16    : inout std_logic := '-';
			wifi_gpio17    : inout std_logic := '-';

			ant_433mhz     : out   std_logic;

			usb_fpga_dp    : inout std_logic := '-';  
			usb_fpga_dn    : inout std_logic := '-';
			usb_fpga_bd_dp : inout std_logic := '-';
			usb_fpga_bd_dn : inout std_logic := '-';
			usb_fpga_pu_dp : inout std_logic := '-';
			usb_fpga_pu_dn : inout std_logic := '-';
						   
			sdram_clk      : inout std_logic;  
			sdram_cke      : out   std_logic;
			sdram_csn      : out   std_logic;
			sdram_wen      : out   std_logic;
			sdram_rasn     : out   std_logic;
			sdram_casn     : out   std_logic;
			sdram_a        : out   std_logic_vector(13-1 downto 0);
			sdram_ba       : out   std_logic_vector(2-1 downto 0);
			sdram_dqm      : inout std_logic_vector(2-1 downto 0) := (others => '-');
			sdram_d        : inout std_logic_vector(16-1 downto 0) := (others => '-');

			gpdi_dp        : out   std_logic_vector(4-1 downto 0);
			gpdi_dn        : out   std_logic_vector(4-1 downto 0);
			--gpdi_ethp      : out   std_logic;  
			--gpdi_ethn      : out   std_logic;
			gpdi_cec       : inout std_logic := '-';
			gpdi_sda       : inout std_logic := '-';
			gpdi_scl       : inout std_logic := '-';

			gp             : inout std_logic_vector(28-1 downto 0) := (others => '-');
			gn             : inout std_logic_vector(28-1 downto 0) := (others => '-');

			user_programn  : out   std_logic := '1'; -- '0' loads next bitstream from SPI FLASH (e.g. bootloader)
			shutdown       : out   std_logic := '0'); -- '1' power off the board, 10uA sleep
	end component;

	component mt48lc32m16a2 is
		port (
			clk   : in std_logic;
			cke   : in std_logic;
			cs_n  : in std_logic;
			ras_n : in std_logic;
			cas_n : in std_logic;
			we_n  : in std_logic;
			ba    : in std_logic_vector(1 downto 0);
			addr  : in std_logic_vector(addr_bits - 1 downto 0);
			dqm   : in std_logic_vector(data_bytes - 1 downto 0);
			dq    : inout std_logic_vector(data_bits - 1 downto 0));
	end component;

	constant baudrate : natural := 115200_00;
	constant uart_data  : std_logic_vector := 
x"000018ff"& 
x"1234ffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffaabb" &
x"ccddffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffff678900001602_5c00_0180_00_00_1702" &
x"5c005c007f000018ffabcdffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffffffff" &
x"ffffffffffffffffffffffffffff50ee" &
x"ffffffffffffffffff00001602_5c00_5c00" &
x"5c00_000017025c005c007f0000";
	
--		x"0000"                             &
--		x"18ff"                             &
--		x"abcd42504250425242924a924a924292" &
--		x"429242524254429442964a966be07420" &
--		x"5b1a5b1a531a531a639e6ba06be06be2" &
--		x"73e274247424742474247c2484aa8cea" &
--		x"84a67c647c647c667c667c24742273e2" &
--		x"7c668cea956e9db0a5b2a5b2a5b2a5b2" &
--		x"a5b09d709d709d709d709db09db09db0" &
--		x"a5b2a5b2a5b2a5b2a5b2a5b2a5f4a5f4" &
--		x"a5f4a5f4adf4adf4adf4adf4adf4adf4" &
--		x"ae34adf4adf4adf4adf4ae34ae34ae34" &
--		x"ae34ae34ae34ae34ae34ae34ae34ae34" &
--		x"ae34ae34ae34ae36b634ae34b634b636" &
--		x"ae34ae34b636b634b636b636b636b636" &
--		x"b634b634b636b636ae34b636b636b636" &
--		x"b634b634b634b634b634b636b636b636" &
--		x"b634b636b636b636b636b636b6364321" &
--		x"0000"                             &
--		x"16025c005c005c00"                 &
--		x"0000"                             &
--		x"17025c005c007f"                   &
--		x"0000"                             &
--		x"18ff"                             &
--		x"1234b636b636b636b636b636b636b636" &
--		x"b636b636b636b636b636b636b636b636" &
--		x"b636b636b636b636b636b636b636b636" &
--		x"b636b636b636b636b636b636b636b636" &
--		x"b636b636b636b636b636b636b636b636" &
--		x"b636b636b636b636b636b636b636b636" &
--		x"b636b636b636b636b636b636b636b636" &
--		x"b636b636b636b636b636b636b636b636" &
--		x"b636b636b636b636b636b636b636b636" &
--		x"b636b636b636b676b676b636b636b636" &
--		x"b676b676b676b676b676b636b636b636" &
--		x"b636b676b676b676b676b676b676b676" &
--		x"b636b676b676b676b676b676b676b636" &
--		x"b676b676b676b676b676b676b676b676" &
--		x"b676b676b676b676b676b676b676be76" &
--		x"b676b676b676b676b676b676b6765a7c" &
--		x"0000"                             &
--		x"16025c005c0080"                   &
--		x"0000"                             &
--		x"17025c005c007f"                   &
--		x"0000";

	signal uart_clk : std_logic := '0';
	signal uart_sin : std_logic;
begin

	rst <= '1', '0' after (1 us+82.5 us);
	xtal <= not xtal after 20 ns;

	uart_clk <= not uart_clk after (1 sec / baudrate / 2);
	process (rst, uart_clk)
		variable data : unsigned((uart_data'length/8)*10-1 downto 0);
	begin
		if rst='1' then
			for i in 0 to data'length/10-1 loop
				data(10-1 downto 0) := unsigned(uart_data(i*8 to (i+1)*8-1)) & b"01";
				data := data ror 10;
			end loop;
			data := not data;
			uart_sin <= '1';
		elsif rising_edge(uart_clk) then
			data := data srl 1;
--			data := data ror 1;
			uart_sin <= not data(0);
		end if;
	end process;

	du_e : ulx3s
	port map (
		clk_25mhz  => xtal,
		ftdi_txd   => uart_sin,

		sdram_clk  => sdram_clk,
		sdram_cke  => sdram_cke,
		sdram_csn  => sdram_cs_n,
		sdram_rasn => sdram_ras_n,
		sdram_casn => sdram_cas_n,
		sdram_wen  => sdram_we_n,
		sdram_ba   => sdram_ba,
		sdram_a    => sdram_addr,
		sdram_dqm  => sdram_dqm,
		sdram_d    => sdram_dq);

	sdr_model_g: mt48lc32m16a2
	port map (
		clk   => sdram_clk,
		cke   => sdram_cke,
		cs_n  => sdram_cs_n,
		ras_n => sdram_ras_n,
		cas_n => sdram_cas_n,
		we_n  => sdram_we_n,
		ba    => sdram_ba,
		addr  => sdram_addr,
		dqm   => sdram_dqm,
		dq    => sdram_dq);
end;

library micron;

configuration ulx3s_structure_md of testbench is
	for ulx3s_graphics
		for all : ulx3s
			use entity work.ulx3s(structure);
		end for;
		for all: mt48lc32m16a2
			use entity micron.mt48lc32m16a2
			port map (
				clk   => sdram_clk,
				cke   => sdram_cke,
				cs_n  => sdram_cs_n,
				ras_n => sdram_ras_n,
				cas_n => sdram_cas_n,
				we_n  => sdram_we_n,
				ba    => sdram_ba,
				addr  => sdram_addr,
				dqm   => sdram_dqm,
				dq    => sdram_dq);
		end for;
	end for;
end;

library micron;

configuration ulx3s_graphics_md of testbench is
	for ulx3s_graphics
		for all : ulx3s
			use entity work.ulx3s(graphics);
		end for;
			for all : mt48lc32m16a2
			use entity micron.mt48lc32m16a2
			port map (
				clk   => sdram_clk,
				cke   => sdram_cke,
				cs_n  => sdram_cs_n,
				ras_n => sdram_ras_n,
				cas_n => sdram_cas_n,
				we_n  => sdram_we_n,
				ba    => sdram_ba,
				addr  => sdram_addr,
				dqm   => sdram_dqm,
				dq    => sdram_dq);
		end for;
	end for;
end;
