library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library unisim;
use unisim.vcomponents.all;

library hdl4fpga;
use hdl4fpga.std.all;

architecture beh of s3estarter is

	constant hz_scales : scale_vector(0 to 16-1) := (
		(from => 0.0, step => 2.50001*5.0*10.0**(-1)),
		(from => 0.0, step => 5.00001*5.0*10.0**(-1)),

		(from => 0.0, step => 1.00001*5.0*10.0**(+0)),
		(from => 0.0, step => 2.50001*5.0*10.0**(+0)),
		(from => 0.0, step => 5.00001*5.0*10.0**(+0)),
                                     
		(from => 0.0, step => 1.00001*5.0*10.0**(+1)),
		(from => 0.0, step => 2.50001*5.0*10.0**(+1)),
		(from => 0.0, step => 5.00001*5.0*10.0**(+1)),
                                     
		(from => 0.0, step => 1.00001*5.0*10.0**(+2)),
		(from => 0.0, step => 2.50001*5.0*10.0**(+2)),
		(from => 0.0, step => 5.00001*5.0*10.0**(+2)),
                                     
		(from => 0.0, step => 1.00001*5.0*10.0**(+3)),
		(from => 0.0, step => 2.50001*5.0*10.0**(+3)),
		(from => 0.0, step => 5.00001*5.0*10.0**(+3)),

		(from => 0.0, step => 1.00001*5.0*10.0**(+4)),
		(from => 0.0, step => 2.50001*5.0*10.0**(+4)));

	constant vt_scales : scale_vector(0 to 16-1) := (
		(from => 7*1.00001*10.0**(+1), step => -1.00001*10.0**(+1)),
		(from => 7*2.50001*10.0**(+1), step => -2.50001*10.0**(+1)),
		(from => 7*5.00001*10.0**(+1), step => -5.00001*10.0**(+1)),

		(from => 7*1.00001*10.0**(-1), step => -1.00001*10.0**(-1)),
		(from => 7*2.50001*10.0**(-1), step => -2.50001*10.0**(-1)),
		(from => 7*5.00001*10.0**(-1), step => -5.00001*10.0**(-1)),

		(from => 7*1.00001*10.0**(+0), step => -1.00001*10.0**(+0)),
		(from => 7*2.50001*10.0**(+0), step => -2.50001*10.0**(+0)),
		(from => 7*5.00001*10.0**(+0), step => -5.00001*10.0**(+0)),

		(from => 7*1.00001*10.0**(+1), step => -1.00001*10.0**(+1)),
		(from => 7*2.50001*10.0**(+1), step => -2.50001*10.0**(+1)),
		(from => 7*5.00001*10.0**(+1), step => -5.00001*10.0**(+1)),

		(from => 7*1.00001*10.0**(-1), step => -1.00001*10.0**(-1)),
		(from => 7*2.50001*10.0**(-1), step => -2.50001*10.0**(-1)),
		(from => 7*5.00001*10.0**(-1), step => -5.00001*10.0**(-1)),

		(from => 7*1.00001*10.0**(+0), step => -1.00001*10.0**(+0)));

	signal sys_clk    : std_logic;
	signal vga_clk    : std_logic;

	constant sample_size : natural := 14;

	function sinctab (
		constant x0 : integer;
		constant x1 : integer;
		constant n  : integer)
		return std_logic_vector is
		variable y   : real;
		variable aux : std_logic_vector(0 to n*(x1-x0+1)-1);
	begin
		for i in 0 to x1-x0 loop
			y := sin(2.0*MATH_PI*real((i+x0))/64.0);
			aux(i*n to (i+1)*n-1) := std_logic_vector(to_unsigned(integer(real(2**(n-2))*y),n));
		end loop;
		return aux;
	end;

	constant inputs : natural := 2;
	signal sample    : std_logic_vector(inputs*sample_size-1 downto 0);
	signal spi_clk   : std_logic;
	signal spiclk_rd : std_logic;
	signal spiclk_fd : std_logic;
	signal sckamp_rd : std_logic;
	signal sckamp_fd : std_logic;
	signal amp_spi   : std_logic;
	signal amp_sdi   : std_logic;
	signal amp_rdy   : std_logic;
	signal adc_spi   : std_logic;
	signal ampcs     : std_logic;
	signal spi_rst   : std_logic;
	signal dac_sdi   : std_logic;
	signal rot_cwse  : std_logic;
	signal rot_rdy   : std_logic;
	signal input_ena : std_logic;
	signal tdiv      : std_logic_vector(4-1 downto 0);
begin

	clkin_ibufg : ibufg
	port map (
		I => xtal,
		O => sys_clk);

	videodcm_e : entity hdl4fpga.dfs
	generic map (
		dcm_per => 20.0,
		dfs_mul => 4,
		dfs_div => 5)
	port map(
		dcm_rst => btn_north,
		dcm_clk => sys_clk,
		dfs_clk => vga_clk);

	spi_b: block
		signal dfs_rst : std_logic;
	begin
		process (btn_north, sys_clk)
			variable cntr : unsigned(0 to 8) := (others => '0');
		begin 
			if btn_north='1' then
				cntr := (others => '0');
			elsif rising_edge(sys_clk) then
				if cntr(0)='0' then
					cntr := cntr + 1;
				end if;
			end if;
			dfs_rst <= not cntr(0);
		end process;

		spidcm_e : entity hdl4fpga.dfs2dfs
		generic map (
			dcm_per  => 20.0,
			dfs1_mul => 32,
			dfs1_div => 25,
			dfs2_mul => 17,
			dfs2_div => 25)
		port map(
			dcm_rst  => dfs_rst,
			dcm_clk  => sys_clk,
			dfs_clk  => spi_clk,
			dcm_lck  => spi_rst);
--		spi_clk <= sys_clk;
--		spi_rst <= not dfs_rst;


		spiclk_rd <= '0' when spi_rst='0' else sckamp_rd when amp_spi='1' else '0' ;
		spiclk_fd <= '0' when spi_rst='0' else sckamp_fd when amp_spi='1' else '1' ;
		spi_mosi  <= amp_sdi   when amp_spi='1' else dac_sdi;

		spi_sck_e : entity hdl4fpga.ddro
		port map (
			clk => spi_clk,
			dr  => spiclk_rd,
			df  => spiclk_fd,
			q   => spi_sck);

		ampclkr_p : process (spi_rst, spi_clk)
			variable cntr : unsigned(0 to 4-1);
		begin
			if spi_rst='0' then
				cntr := (others => '0');
				sckamp_rd <= cntr(0);
				adc_spi <= '1';
			elsif rising_edge(spi_clk) then
				cntr := cntr + 1;
				sckamp_rd <= cntr(0);
				amp_cs <= ampcs;
			end if;
		end process;

		ampclkf_p : process (spi_rst, spi_clk)
		begin
			if spi_rst='0' then
				sckamp_fd <= '0';
			elsif falling_edge(spi_clk) then
				sckamp_fd <= sckamp_rd;
			end if;
		end process;

		ampp2sr_p : process (spi_rst, sckamp_fd)
		begin
			if spi_rst='0' then
				ampcs <= '1';
			elsif falling_edge(sckamp_fd) then
				ampcs <= not amp_rdy or not amp_spi;
			end if;
		end process;

		amp_p : process (spi_rst, sckamp_fd)
			variable cntr : unsigned(0 to 4);
			variable val  : unsigned(0 to 8-1);
		begin
			if spi_rst='0' then
				amp_spi <= '1';
				amp_rdy <= '0';
				amp_sdi <= '0';
				cntr    := to_unsigned(val'length-2,cntr'length);
				val     := B"0001_0001";
			elsif falling_edge(sckamp_fd) then
				if ampcs='0' then
					if cntr(0)='0' then
						cntr := cntr - 1;
						val  := val rol 1;
					end if;
				end if;
				amp_sdi <= val(0);
				amp_rdy <= not cntr(0);
				amp_spi <= not cntr(0) or not ampcs;
			end if;
		end process;

		adcdac_p : process (amp_spi, spi_clk)
			constant p2p        : natural := 2*1550;
			constant cycle      : natural := 34;
			variable cntr       : unsigned(0 to 6) := (others => '0');
			variable adin       : unsigned(32-1 downto 0);
			variable aux        : unsigned(sample'range);
			variable dac_shr    : unsigned(0 to 30-1);
			variable adcdac_sel : std_logic;
			variable dac_data   : unsigned(0 to 12-1);
			variable dac_chan   : unsigned(0 to 2-1);
		begin
			if amp_spi='1' then
				cntr       := to_unsigned(cycle-2, cntr'length);
				adcdac_sel := '0';
				dac_sdi    <= '0';
				dac_cs     <= '1';
			elsif rising_edge(spi_clk) then
				if cntr(0)='1' then
					if adcdac_sel ='0' then

--						for i in 0 to inputs-1 loop
--							aux := aux sll sample_size;
--							aux(sample_size-1 downto 0) := not adin(sample_size-1 downto 0);
--							adin := adin srl (adin'length/inputs);
--						end loop;
--						sample <= std_logic_vector(aux);
						sample <= std_logic_vector(
							not adin(1*16+sample_size-1 downto 1*16) &
							not adin(0*16+sample_size-1 downto 0*16));

						input_ena <= not amp_spi;
						ad_conv   <= '0';
					else
						if to_integer(dac_data)=(2048+p2p/2) then
							dac_data := to_unsigned(2048-p2p/2, dac_data'length);
						else
							dac_data := dac_data + 1;
						end if;
						ad_conv <= not amp_spi;
					end if;

					if tdiv=(1 to 4 => '0') then
						adcdac_sel := '0';
						ad_conv    <= '1';
					else 
						adcdac_sel := not adcdac_sel;
					end if;

					dac_shr := (1 to 10 => '-') & "001100" & dac_chan & dac_data;
					cntr    := to_unsigned(cycle-2, cntr'length);
				else
					input_ena <= '0';
					ad_conv   <= '0';
					dac_shr   := dac_shr sll 1;
					cntr      := cntr - 1;
				end if;
				adin    := adin sll 1;
				adin(0) := spi_miso;

				dac_cs  <= not adcdac_sel or amp_spi;
				dac_sdi <= dac_shr(0);
			end if;
		end process;
	end block;

	process (e_rx_clk, rot_a, rot_b)
		variable cntr : unsigned(0 to 12);
	begin
		if (rot_a or rot_b)='1' then
			if cntr(0)='1' then
				cntr := (others => '0');
			end if;
			rot_cwse <= rot_a;
		elsif rising_edge(xtal) then
			if cntr(0)='0' then
				cntr := cntr + 1;
			end if;
			rot_rdy <= cntr(0);
		end if;
	end process;

	scopeio_e : entity hdl4fpga.scopeio
	generic map (
		layout_id  => 1,
		hz_scales  => hz_scales,
		vt_scales  => vt_scales,
		inputs => inputs,
		input_unit => 100.0*(1.25*64.0)/8192.0)
	port map (
		mii_rxc     => e_rx_clk,
		mii_rxdv    => e_rx_dv,
		mii_rxd     => e_rxd,
		tdiv        => tdiv,
		input_clk   => spi_clk,
		input_ena   => input_ena,
		input_data  => sample,
		video_clk   => vga_clk,
		video_red   => vga_red,
		video_green => vga_green,
		video_blue  => vga_blue,
		video_hsync => vga_hsync,
		video_vsync => vga_vsync);

	-- Ethernet Transceiver --
	--------------------------

	e_txen <= 'Z';
	e_txd  <= (others => 'Z');
	e_mdc  <= '0';
	e_mdio <= 'Z';
	e_txd_4 <= '0';

	-- DDR --
	---------

	ddr_clk_i : obufds
	generic map (
		iostandard => "DIFF_SSTL2_I")
	port map (
		i  => 'Z',
		o  => sd_ck_p,
		ob => sd_ck_n);

	sd_cke    <= 'Z';
	sd_cs     <= 'Z';
	sd_ras    <= 'Z';
	sd_cas    <= 'Z';
	sd_we     <= 'Z';
	sd_ba     <= (others => 'Z');
	sd_a      <= (others => 'Z');
	sd_dm     <= (others => 'Z');
	sd_dqs    <= (others => 'Z');
	sd_dq     <= (others => 'Z');

	amp_shdn <= '0';
	dac_clr <= '1';
	sf_ce0 <= '1';
	fpga_init_b <= '0';
	spi_ss_b <= '0';

	led0 <= '1';
	led1 <= '1';
	led2 <= '1';
	led3 <= '1';
	led4 <= '1';
	led5 <= '1';
	led6 <= '1';
	led7 <= '1';
end;
