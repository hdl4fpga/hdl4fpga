constant psf1unitx8x8 : std_logic_vector(0 to 16*8*8-1) := (
	"01111100" &
	"11001110" &
	"11011110" &
	"11110110" &
	"11100110" &
	"11000110" &
	"01111100" &
	"00000000" &

	"00011000" &
	"00111000" &
	"00011000" &
	"00011000" &
	"00011000" &
	"00011000" &
	"01111110" &
	"00000000" &

	"01111100" &
	"11000110" &
	"00000110" &
	"01111100" &
	"11000000" &
	"11000000" &
	"11111110" &
	"00000000" &

	"11111100" &
	"00000110" &
	"00000110" &
	"00111100" &
	"00000110" &
	"00000110" &
	"11111100" &
	"00000000" &

	"00001100" &
	"11001100" &
	"11001100" &
	"11001100" &
	"11111110" &
	"00001100" &
	"00001100" &
	"00000000" &

	"11111110" &
	"11000000" &
	"11111100" &
	"00000110" &
	"00000110" &
	"11000110" &
	"01111100" &
	"00000000" &

	"01111100" &
	"11000000" &
	"11000000" &
	"11111100" &
	"11000110" &
	"11000110" &
	"01111100" &
	"00000000" &

	"11111110" &
	"00000110" &
	"00000110" &
	"00001100" &
	"00011000" &
	"00110000" &
	"00110000" &
	"00000000" &

	"01111100" &
	"11000110" &
	"11000110" &
	"01111100" &
	"11000110" &
	"11000110" &
	"01111100" &
	"00000000" &

	"01111100" &
	"11000110" &
	"11000110" &
	"01111110" &
	"00000110" &
	"00000110" &
	"01111100" &
	"00000000" &

	"00000000" &
	"00000000" &
	"00000000" &
	"00000000" &
	"00000000" &
	"00011000" &
	"00011000" &
	"00000000" &

	"00000000" &
	"00000000" &
	"11001100" &
	"11111110" &
	"11111110" &
	"11010110" &
	"11010110" &
	"00000000" &

	"00000000" &
	"00000000" &
	"11111100" &
	"11000110" &
	"11000110" &
	"11000110" &
	"11000110" &
	"00000000" &

	"00000000" &
	"01100110" &
	"01100110" &
	"01100110" &
	"01100110" &
	"01111100" &
	"01100000" &
	"11000000");

	"11000110" &
	"11000110" &
	"11000110" &
	"11000110" &
	"11000110" &
	"01111100" &
	"00111000" &
	"00000000" &

	"00000000" &
	"00000000" &
	"01111110" &
	"11000000" &
	"01111100" &
	"00000110" &
	"11111100" &
	"00000000");
